magic
tech sky130A
magscale 1 2
timestamp 1717069679
<< viali >>
rect 7021 6817 7055 6851
rect 6837 6613 6871 6647
rect 3433 6341 3467 6375
rect 3985 6205 4019 6239
rect 4445 6205 4479 6239
rect 4997 6205 5031 6239
rect 5549 6205 5583 6239
rect 3801 6137 3835 6171
rect 3341 6069 3375 6103
rect 4077 6069 4111 6103
rect 4353 6069 4387 6103
rect 2421 5797 2455 5831
rect 2789 5797 2823 5831
rect 2973 5797 3007 5831
rect 4077 5797 4111 5831
rect 3249 5729 3283 5763
rect 3709 5729 3743 5763
rect 3801 5729 3835 5763
rect 5549 5661 5583 5695
rect 3709 5321 3743 5355
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
<< metal1 >>
rect 552 7098 7520 7120
rect 552 7046 2100 7098
rect 2152 7046 2164 7098
rect 2216 7046 2228 7098
rect 2280 7046 2292 7098
rect 2344 7046 2356 7098
rect 2408 7046 3802 7098
rect 3854 7046 3866 7098
rect 3918 7046 3930 7098
rect 3982 7046 3994 7098
rect 4046 7046 4058 7098
rect 4110 7046 5504 7098
rect 5556 7046 5568 7098
rect 5620 7046 5632 7098
rect 5684 7046 5696 7098
rect 5748 7046 5760 7098
rect 5812 7046 7206 7098
rect 7258 7046 7270 7098
rect 7322 7046 7334 7098
rect 7386 7046 7398 7098
rect 7450 7046 7462 7098
rect 7514 7046 7520 7098
rect 552 7024 7520 7046
rect 6822 6944 6828 6996
rect 6880 6944 6886 6996
rect 6840 6848 6868 6944
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6840 6820 7021 6848
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 5408 6616 6837 6644
rect 5408 6604 5414 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 552 6554 7360 6576
rect 552 6502 1249 6554
rect 1301 6502 1313 6554
rect 1365 6502 1377 6554
rect 1429 6502 1441 6554
rect 1493 6502 1505 6554
rect 1557 6502 2951 6554
rect 3003 6502 3015 6554
rect 3067 6502 3079 6554
rect 3131 6502 3143 6554
rect 3195 6502 3207 6554
rect 3259 6502 4653 6554
rect 4705 6502 4717 6554
rect 4769 6502 4781 6554
rect 4833 6502 4845 6554
rect 4897 6502 4909 6554
rect 4961 6502 6355 6554
rect 6407 6502 6419 6554
rect 6471 6502 6483 6554
rect 6535 6502 6547 6554
rect 6599 6502 6611 6554
rect 6663 6502 7360 6554
rect 552 6480 7360 6502
rect 3418 6332 3424 6384
rect 3476 6332 3482 6384
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4479 6208 4997 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 3789 6171 3847 6177
rect 3789 6168 3801 6171
rect 3752 6140 3801 6168
rect 3752 6128 3758 6140
rect 3789 6137 3801 6140
rect 3835 6168 3847 6171
rect 3988 6168 4016 6199
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5316 6208 5549 6236
rect 5316 6196 5322 6208
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 3835 6140 4016 6168
rect 3835 6137 3847 6140
rect 3789 6131 3847 6137
rect 3326 6060 3332 6112
rect 3384 6060 3390 6112
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4154 6100 4160 6112
rect 4111 6072 4160 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 4338 6060 4344 6112
rect 4396 6060 4402 6112
rect 552 6010 7520 6032
rect 552 5958 2100 6010
rect 2152 5958 2164 6010
rect 2216 5958 2228 6010
rect 2280 5958 2292 6010
rect 2344 5958 2356 6010
rect 2408 5958 3802 6010
rect 3854 5958 3866 6010
rect 3918 5958 3930 6010
rect 3982 5958 3994 6010
rect 4046 5958 4058 6010
rect 4110 5958 5504 6010
rect 5556 5958 5568 6010
rect 5620 5958 5632 6010
rect 5684 5958 5696 6010
rect 5748 5958 5760 6010
rect 5812 5958 7206 6010
rect 7258 5958 7270 6010
rect 7322 5958 7334 6010
rect 7386 5958 7398 6010
rect 7450 5958 7462 6010
rect 7514 5958 7520 6010
rect 552 5936 7520 5958
rect 3326 5896 3332 5908
rect 2792 5868 3332 5896
rect 1578 5788 1584 5840
rect 1636 5828 1642 5840
rect 2792 5837 2820 5868
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 4982 5896 4988 5908
rect 3804 5868 4988 5896
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 1636 5800 2421 5828
rect 1636 5788 1642 5800
rect 2409 5797 2421 5800
rect 2455 5797 2467 5831
rect 2409 5791 2467 5797
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5797 2835 5831
rect 2777 5791 2835 5797
rect 2958 5788 2964 5840
rect 3016 5788 3022 5840
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 3436 5760 3464 5856
rect 3283 5732 3464 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 3436 5692 3464 5732
rect 3694 5720 3700 5772
rect 3752 5720 3758 5772
rect 3804 5769 3832 5868
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 4065 5831 4123 5837
rect 4065 5797 4077 5831
rect 4111 5828 4123 5831
rect 4338 5828 4344 5840
rect 4111 5800 4344 5828
rect 4111 5797 4123 5800
rect 4065 5791 4123 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5350 5828 5356 5840
rect 5290 5800 5356 5828
rect 5350 5788 5356 5800
rect 5408 5788 5414 5840
rect 3789 5763 3847 5769
rect 3789 5729 3801 5763
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 5258 5692 5264 5704
rect 3436 5664 5264 5692
rect 5258 5652 5264 5664
rect 5316 5692 5322 5704
rect 5442 5692 5448 5704
rect 5316 5664 5448 5692
rect 5316 5652 5322 5664
rect 5442 5652 5448 5664
rect 5500 5692 5506 5704
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5500 5664 5549 5692
rect 5500 5652 5506 5664
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 552 5466 7360 5488
rect 552 5414 1249 5466
rect 1301 5414 1313 5466
rect 1365 5414 1377 5466
rect 1429 5414 1441 5466
rect 1493 5414 1505 5466
rect 1557 5414 2951 5466
rect 3003 5414 3015 5466
rect 3067 5414 3079 5466
rect 3131 5414 3143 5466
rect 3195 5414 3207 5466
rect 3259 5414 4653 5466
rect 4705 5414 4717 5466
rect 4769 5414 4781 5466
rect 4833 5414 4845 5466
rect 4897 5414 4909 5466
rect 4961 5414 6355 5466
rect 6407 5414 6419 5466
rect 6471 5414 6483 5466
rect 6535 5414 6547 5466
rect 6599 5414 6611 5466
rect 6663 5414 7360 5466
rect 552 5392 7360 5414
rect 3694 5312 3700 5364
rect 3752 5312 3758 5364
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 4172 5216 4200 5312
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4172 5188 5181 5216
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 4738 5052 5396 5080
rect 5368 5024 5396 5052
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 552 4922 7520 4944
rect 552 4870 2100 4922
rect 2152 4870 2164 4922
rect 2216 4870 2228 4922
rect 2280 4870 2292 4922
rect 2344 4870 2356 4922
rect 2408 4870 3802 4922
rect 3854 4870 3866 4922
rect 3918 4870 3930 4922
rect 3982 4870 3994 4922
rect 4046 4870 4058 4922
rect 4110 4870 5504 4922
rect 5556 4870 5568 4922
rect 5620 4870 5632 4922
rect 5684 4870 5696 4922
rect 5748 4870 5760 4922
rect 5812 4870 7206 4922
rect 7258 4870 7270 4922
rect 7322 4870 7334 4922
rect 7386 4870 7398 4922
rect 7450 4870 7462 4922
rect 7514 4870 7520 4922
rect 552 4848 7520 4870
rect 552 4378 7360 4400
rect 552 4326 1249 4378
rect 1301 4326 1313 4378
rect 1365 4326 1377 4378
rect 1429 4326 1441 4378
rect 1493 4326 1505 4378
rect 1557 4326 2951 4378
rect 3003 4326 3015 4378
rect 3067 4326 3079 4378
rect 3131 4326 3143 4378
rect 3195 4326 3207 4378
rect 3259 4326 4653 4378
rect 4705 4326 4717 4378
rect 4769 4326 4781 4378
rect 4833 4326 4845 4378
rect 4897 4326 4909 4378
rect 4961 4326 6355 4378
rect 6407 4326 6419 4378
rect 6471 4326 6483 4378
rect 6535 4326 6547 4378
rect 6599 4326 6611 4378
rect 6663 4326 7360 4378
rect 552 4304 7360 4326
rect 552 3834 7520 3856
rect 552 3782 2100 3834
rect 2152 3782 2164 3834
rect 2216 3782 2228 3834
rect 2280 3782 2292 3834
rect 2344 3782 2356 3834
rect 2408 3782 3802 3834
rect 3854 3782 3866 3834
rect 3918 3782 3930 3834
rect 3982 3782 3994 3834
rect 4046 3782 4058 3834
rect 4110 3782 5504 3834
rect 5556 3782 5568 3834
rect 5620 3782 5632 3834
rect 5684 3782 5696 3834
rect 5748 3782 5760 3834
rect 5812 3782 7206 3834
rect 7258 3782 7270 3834
rect 7322 3782 7334 3834
rect 7386 3782 7398 3834
rect 7450 3782 7462 3834
rect 7514 3782 7520 3834
rect 552 3760 7520 3782
rect 552 3290 7360 3312
rect 552 3238 1249 3290
rect 1301 3238 1313 3290
rect 1365 3238 1377 3290
rect 1429 3238 1441 3290
rect 1493 3238 1505 3290
rect 1557 3238 2951 3290
rect 3003 3238 3015 3290
rect 3067 3238 3079 3290
rect 3131 3238 3143 3290
rect 3195 3238 3207 3290
rect 3259 3238 4653 3290
rect 4705 3238 4717 3290
rect 4769 3238 4781 3290
rect 4833 3238 4845 3290
rect 4897 3238 4909 3290
rect 4961 3238 6355 3290
rect 6407 3238 6419 3290
rect 6471 3238 6483 3290
rect 6535 3238 6547 3290
rect 6599 3238 6611 3290
rect 6663 3238 7360 3290
rect 552 3216 7360 3238
rect 552 2746 7520 2768
rect 552 2694 2100 2746
rect 2152 2694 2164 2746
rect 2216 2694 2228 2746
rect 2280 2694 2292 2746
rect 2344 2694 2356 2746
rect 2408 2694 3802 2746
rect 3854 2694 3866 2746
rect 3918 2694 3930 2746
rect 3982 2694 3994 2746
rect 4046 2694 4058 2746
rect 4110 2694 5504 2746
rect 5556 2694 5568 2746
rect 5620 2694 5632 2746
rect 5684 2694 5696 2746
rect 5748 2694 5760 2746
rect 5812 2694 7206 2746
rect 7258 2694 7270 2746
rect 7322 2694 7334 2746
rect 7386 2694 7398 2746
rect 7450 2694 7462 2746
rect 7514 2694 7520 2746
rect 552 2672 7520 2694
rect 552 2202 7360 2224
rect 552 2150 1249 2202
rect 1301 2150 1313 2202
rect 1365 2150 1377 2202
rect 1429 2150 1441 2202
rect 1493 2150 1505 2202
rect 1557 2150 2951 2202
rect 3003 2150 3015 2202
rect 3067 2150 3079 2202
rect 3131 2150 3143 2202
rect 3195 2150 3207 2202
rect 3259 2150 4653 2202
rect 4705 2150 4717 2202
rect 4769 2150 4781 2202
rect 4833 2150 4845 2202
rect 4897 2150 4909 2202
rect 4961 2150 6355 2202
rect 6407 2150 6419 2202
rect 6471 2150 6483 2202
rect 6535 2150 6547 2202
rect 6599 2150 6611 2202
rect 6663 2150 7360 2202
rect 552 2128 7360 2150
rect 552 1658 7520 1680
rect 552 1606 2100 1658
rect 2152 1606 2164 1658
rect 2216 1606 2228 1658
rect 2280 1606 2292 1658
rect 2344 1606 2356 1658
rect 2408 1606 3802 1658
rect 3854 1606 3866 1658
rect 3918 1606 3930 1658
rect 3982 1606 3994 1658
rect 4046 1606 4058 1658
rect 4110 1606 5504 1658
rect 5556 1606 5568 1658
rect 5620 1606 5632 1658
rect 5684 1606 5696 1658
rect 5748 1606 5760 1658
rect 5812 1606 7206 1658
rect 7258 1606 7270 1658
rect 7322 1606 7334 1658
rect 7386 1606 7398 1658
rect 7450 1606 7462 1658
rect 7514 1606 7520 1658
rect 552 1584 7520 1606
rect 552 1114 7360 1136
rect 552 1062 1249 1114
rect 1301 1062 1313 1114
rect 1365 1062 1377 1114
rect 1429 1062 1441 1114
rect 1493 1062 1505 1114
rect 1557 1062 2951 1114
rect 3003 1062 3015 1114
rect 3067 1062 3079 1114
rect 3131 1062 3143 1114
rect 3195 1062 3207 1114
rect 3259 1062 4653 1114
rect 4705 1062 4717 1114
rect 4769 1062 4781 1114
rect 4833 1062 4845 1114
rect 4897 1062 4909 1114
rect 4961 1062 6355 1114
rect 6407 1062 6419 1114
rect 6471 1062 6483 1114
rect 6535 1062 6547 1114
rect 6599 1062 6611 1114
rect 6663 1062 7360 1114
rect 552 1040 7360 1062
rect 552 570 7520 592
rect 552 518 2100 570
rect 2152 518 2164 570
rect 2216 518 2228 570
rect 2280 518 2292 570
rect 2344 518 2356 570
rect 2408 518 3802 570
rect 3854 518 3866 570
rect 3918 518 3930 570
rect 3982 518 3994 570
rect 4046 518 4058 570
rect 4110 518 5504 570
rect 5556 518 5568 570
rect 5620 518 5632 570
rect 5684 518 5696 570
rect 5748 518 5760 570
rect 5812 518 7206 570
rect 7258 518 7270 570
rect 7322 518 7334 570
rect 7386 518 7398 570
rect 7450 518 7462 570
rect 7514 518 7520 570
rect 552 496 7520 518
<< via1 >>
rect 2100 7046 2152 7098
rect 2164 7046 2216 7098
rect 2228 7046 2280 7098
rect 2292 7046 2344 7098
rect 2356 7046 2408 7098
rect 3802 7046 3854 7098
rect 3866 7046 3918 7098
rect 3930 7046 3982 7098
rect 3994 7046 4046 7098
rect 4058 7046 4110 7098
rect 5504 7046 5556 7098
rect 5568 7046 5620 7098
rect 5632 7046 5684 7098
rect 5696 7046 5748 7098
rect 5760 7046 5812 7098
rect 7206 7046 7258 7098
rect 7270 7046 7322 7098
rect 7334 7046 7386 7098
rect 7398 7046 7450 7098
rect 7462 7046 7514 7098
rect 6828 6944 6880 6996
rect 5356 6604 5408 6656
rect 1249 6502 1301 6554
rect 1313 6502 1365 6554
rect 1377 6502 1429 6554
rect 1441 6502 1493 6554
rect 1505 6502 1557 6554
rect 2951 6502 3003 6554
rect 3015 6502 3067 6554
rect 3079 6502 3131 6554
rect 3143 6502 3195 6554
rect 3207 6502 3259 6554
rect 4653 6502 4705 6554
rect 4717 6502 4769 6554
rect 4781 6502 4833 6554
rect 4845 6502 4897 6554
rect 4909 6502 4961 6554
rect 6355 6502 6407 6554
rect 6419 6502 6471 6554
rect 6483 6502 6535 6554
rect 6547 6502 6599 6554
rect 6611 6502 6663 6554
rect 3424 6375 3476 6384
rect 3424 6341 3433 6375
rect 3433 6341 3467 6375
rect 3467 6341 3476 6375
rect 3424 6332 3476 6341
rect 3700 6128 3752 6180
rect 5264 6196 5316 6248
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 4160 6060 4212 6112
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 2100 5958 2152 6010
rect 2164 5958 2216 6010
rect 2228 5958 2280 6010
rect 2292 5958 2344 6010
rect 2356 5958 2408 6010
rect 3802 5958 3854 6010
rect 3866 5958 3918 6010
rect 3930 5958 3982 6010
rect 3994 5958 4046 6010
rect 4058 5958 4110 6010
rect 5504 5958 5556 6010
rect 5568 5958 5620 6010
rect 5632 5958 5684 6010
rect 5696 5958 5748 6010
rect 5760 5958 5812 6010
rect 7206 5958 7258 6010
rect 7270 5958 7322 6010
rect 7334 5958 7386 6010
rect 7398 5958 7450 6010
rect 7462 5958 7514 6010
rect 1584 5788 1636 5840
rect 3332 5856 3384 5908
rect 3424 5856 3476 5908
rect 2964 5831 3016 5840
rect 2964 5797 2973 5831
rect 2973 5797 3007 5831
rect 3007 5797 3016 5831
rect 2964 5788 3016 5797
rect 3700 5763 3752 5772
rect 3700 5729 3709 5763
rect 3709 5729 3743 5763
rect 3743 5729 3752 5763
rect 3700 5720 3752 5729
rect 4988 5856 5040 5908
rect 4344 5788 4396 5840
rect 5356 5788 5408 5840
rect 5264 5652 5316 5704
rect 5448 5652 5500 5704
rect 1249 5414 1301 5466
rect 1313 5414 1365 5466
rect 1377 5414 1429 5466
rect 1441 5414 1493 5466
rect 1505 5414 1557 5466
rect 2951 5414 3003 5466
rect 3015 5414 3067 5466
rect 3079 5414 3131 5466
rect 3143 5414 3195 5466
rect 3207 5414 3259 5466
rect 4653 5414 4705 5466
rect 4717 5414 4769 5466
rect 4781 5414 4833 5466
rect 4845 5414 4897 5466
rect 4909 5414 4961 5466
rect 6355 5414 6407 5466
rect 6419 5414 6471 5466
rect 6483 5414 6535 5466
rect 6547 5414 6599 5466
rect 6611 5414 6663 5466
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 4160 5312 4212 5364
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 5356 4972 5408 5024
rect 2100 4870 2152 4922
rect 2164 4870 2216 4922
rect 2228 4870 2280 4922
rect 2292 4870 2344 4922
rect 2356 4870 2408 4922
rect 3802 4870 3854 4922
rect 3866 4870 3918 4922
rect 3930 4870 3982 4922
rect 3994 4870 4046 4922
rect 4058 4870 4110 4922
rect 5504 4870 5556 4922
rect 5568 4870 5620 4922
rect 5632 4870 5684 4922
rect 5696 4870 5748 4922
rect 5760 4870 5812 4922
rect 7206 4870 7258 4922
rect 7270 4870 7322 4922
rect 7334 4870 7386 4922
rect 7398 4870 7450 4922
rect 7462 4870 7514 4922
rect 1249 4326 1301 4378
rect 1313 4326 1365 4378
rect 1377 4326 1429 4378
rect 1441 4326 1493 4378
rect 1505 4326 1557 4378
rect 2951 4326 3003 4378
rect 3015 4326 3067 4378
rect 3079 4326 3131 4378
rect 3143 4326 3195 4378
rect 3207 4326 3259 4378
rect 4653 4326 4705 4378
rect 4717 4326 4769 4378
rect 4781 4326 4833 4378
rect 4845 4326 4897 4378
rect 4909 4326 4961 4378
rect 6355 4326 6407 4378
rect 6419 4326 6471 4378
rect 6483 4326 6535 4378
rect 6547 4326 6599 4378
rect 6611 4326 6663 4378
rect 2100 3782 2152 3834
rect 2164 3782 2216 3834
rect 2228 3782 2280 3834
rect 2292 3782 2344 3834
rect 2356 3782 2408 3834
rect 3802 3782 3854 3834
rect 3866 3782 3918 3834
rect 3930 3782 3982 3834
rect 3994 3782 4046 3834
rect 4058 3782 4110 3834
rect 5504 3782 5556 3834
rect 5568 3782 5620 3834
rect 5632 3782 5684 3834
rect 5696 3782 5748 3834
rect 5760 3782 5812 3834
rect 7206 3782 7258 3834
rect 7270 3782 7322 3834
rect 7334 3782 7386 3834
rect 7398 3782 7450 3834
rect 7462 3782 7514 3834
rect 1249 3238 1301 3290
rect 1313 3238 1365 3290
rect 1377 3238 1429 3290
rect 1441 3238 1493 3290
rect 1505 3238 1557 3290
rect 2951 3238 3003 3290
rect 3015 3238 3067 3290
rect 3079 3238 3131 3290
rect 3143 3238 3195 3290
rect 3207 3238 3259 3290
rect 4653 3238 4705 3290
rect 4717 3238 4769 3290
rect 4781 3238 4833 3290
rect 4845 3238 4897 3290
rect 4909 3238 4961 3290
rect 6355 3238 6407 3290
rect 6419 3238 6471 3290
rect 6483 3238 6535 3290
rect 6547 3238 6599 3290
rect 6611 3238 6663 3290
rect 2100 2694 2152 2746
rect 2164 2694 2216 2746
rect 2228 2694 2280 2746
rect 2292 2694 2344 2746
rect 2356 2694 2408 2746
rect 3802 2694 3854 2746
rect 3866 2694 3918 2746
rect 3930 2694 3982 2746
rect 3994 2694 4046 2746
rect 4058 2694 4110 2746
rect 5504 2694 5556 2746
rect 5568 2694 5620 2746
rect 5632 2694 5684 2746
rect 5696 2694 5748 2746
rect 5760 2694 5812 2746
rect 7206 2694 7258 2746
rect 7270 2694 7322 2746
rect 7334 2694 7386 2746
rect 7398 2694 7450 2746
rect 7462 2694 7514 2746
rect 1249 2150 1301 2202
rect 1313 2150 1365 2202
rect 1377 2150 1429 2202
rect 1441 2150 1493 2202
rect 1505 2150 1557 2202
rect 2951 2150 3003 2202
rect 3015 2150 3067 2202
rect 3079 2150 3131 2202
rect 3143 2150 3195 2202
rect 3207 2150 3259 2202
rect 4653 2150 4705 2202
rect 4717 2150 4769 2202
rect 4781 2150 4833 2202
rect 4845 2150 4897 2202
rect 4909 2150 4961 2202
rect 6355 2150 6407 2202
rect 6419 2150 6471 2202
rect 6483 2150 6535 2202
rect 6547 2150 6599 2202
rect 6611 2150 6663 2202
rect 2100 1606 2152 1658
rect 2164 1606 2216 1658
rect 2228 1606 2280 1658
rect 2292 1606 2344 1658
rect 2356 1606 2408 1658
rect 3802 1606 3854 1658
rect 3866 1606 3918 1658
rect 3930 1606 3982 1658
rect 3994 1606 4046 1658
rect 4058 1606 4110 1658
rect 5504 1606 5556 1658
rect 5568 1606 5620 1658
rect 5632 1606 5684 1658
rect 5696 1606 5748 1658
rect 5760 1606 5812 1658
rect 7206 1606 7258 1658
rect 7270 1606 7322 1658
rect 7334 1606 7386 1658
rect 7398 1606 7450 1658
rect 7462 1606 7514 1658
rect 1249 1062 1301 1114
rect 1313 1062 1365 1114
rect 1377 1062 1429 1114
rect 1441 1062 1493 1114
rect 1505 1062 1557 1114
rect 2951 1062 3003 1114
rect 3015 1062 3067 1114
rect 3079 1062 3131 1114
rect 3143 1062 3195 1114
rect 3207 1062 3259 1114
rect 4653 1062 4705 1114
rect 4717 1062 4769 1114
rect 4781 1062 4833 1114
rect 4845 1062 4897 1114
rect 4909 1062 4961 1114
rect 6355 1062 6407 1114
rect 6419 1062 6471 1114
rect 6483 1062 6535 1114
rect 6547 1062 6599 1114
rect 6611 1062 6663 1114
rect 2100 518 2152 570
rect 2164 518 2216 570
rect 2228 518 2280 570
rect 2292 518 2344 570
rect 2356 518 2408 570
rect 3802 518 3854 570
rect 3866 518 3918 570
rect 3930 518 3982 570
rect 3994 518 4046 570
rect 4058 518 4110 570
rect 5504 518 5556 570
rect 5568 518 5620 570
rect 5632 518 5684 570
rect 5696 518 5748 570
rect 5760 518 5812 570
rect 7206 518 7258 570
rect 7270 518 7322 570
rect 7334 518 7386 570
rect 7398 518 7450 570
rect 7462 518 7514 570
<< metal2 >>
rect 1030 7698 1086 8000
rect 2962 7698 3018 8000
rect 1030 7670 1624 7698
rect 1030 7600 1086 7670
rect 1249 6556 1557 6565
rect 1249 6554 1255 6556
rect 1311 6554 1335 6556
rect 1391 6554 1415 6556
rect 1471 6554 1495 6556
rect 1551 6554 1557 6556
rect 1311 6502 1313 6554
rect 1493 6502 1495 6554
rect 1249 6500 1255 6502
rect 1311 6500 1335 6502
rect 1391 6500 1415 6502
rect 1471 6500 1495 6502
rect 1551 6500 1557 6502
rect 1249 6491 1557 6500
rect 1596 5846 1624 7670
rect 2884 7670 3018 7698
rect 2100 7100 2408 7109
rect 2100 7098 2106 7100
rect 2162 7098 2186 7100
rect 2242 7098 2266 7100
rect 2322 7098 2346 7100
rect 2402 7098 2408 7100
rect 2162 7046 2164 7098
rect 2344 7046 2346 7098
rect 2100 7044 2106 7046
rect 2162 7044 2186 7046
rect 2242 7044 2266 7046
rect 2322 7044 2346 7046
rect 2402 7044 2408 7046
rect 2100 7035 2408 7044
rect 2884 6338 2912 7670
rect 2962 7600 3018 7670
rect 4894 7698 4950 8000
rect 4894 7670 5028 7698
rect 4894 7600 4950 7670
rect 3802 7100 4110 7109
rect 3802 7098 3808 7100
rect 3864 7098 3888 7100
rect 3944 7098 3968 7100
rect 4024 7098 4048 7100
rect 4104 7098 4110 7100
rect 3864 7046 3866 7098
rect 4046 7046 4048 7098
rect 3802 7044 3808 7046
rect 3864 7044 3888 7046
rect 3944 7044 3968 7046
rect 4024 7044 4048 7046
rect 4104 7044 4110 7046
rect 3802 7035 4110 7044
rect 2951 6556 3259 6565
rect 2951 6554 2957 6556
rect 3013 6554 3037 6556
rect 3093 6554 3117 6556
rect 3173 6554 3197 6556
rect 3253 6554 3259 6556
rect 3013 6502 3015 6554
rect 3195 6502 3197 6554
rect 2951 6500 2957 6502
rect 3013 6500 3037 6502
rect 3093 6500 3117 6502
rect 3173 6500 3197 6502
rect 3253 6500 3259 6502
rect 2951 6491 3259 6500
rect 4653 6556 4961 6565
rect 4653 6554 4659 6556
rect 4715 6554 4739 6556
rect 4795 6554 4819 6556
rect 4875 6554 4899 6556
rect 4955 6554 4961 6556
rect 4715 6502 4717 6554
rect 4897 6502 4899 6554
rect 4653 6500 4659 6502
rect 4715 6500 4739 6502
rect 4795 6500 4819 6502
rect 4875 6500 4899 6502
rect 4955 6500 4961 6502
rect 4653 6491 4961 6500
rect 3424 6384 3476 6390
rect 2884 6310 3004 6338
rect 3424 6326 3476 6332
rect 2100 6012 2408 6021
rect 2100 6010 2106 6012
rect 2162 6010 2186 6012
rect 2242 6010 2266 6012
rect 2322 6010 2346 6012
rect 2402 6010 2408 6012
rect 2162 5958 2164 6010
rect 2344 5958 2346 6010
rect 2100 5956 2106 5958
rect 2162 5956 2186 5958
rect 2242 5956 2266 5958
rect 2322 5956 2346 5958
rect 2402 5956 2408 5958
rect 2100 5947 2408 5956
rect 2976 5846 3004 6310
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5914 3372 6054
rect 3436 5914 3464 6326
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 1584 5840 1636 5846
rect 1584 5782 1636 5788
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 3712 5778 3740 6122
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 3802 6012 4110 6021
rect 3802 6010 3808 6012
rect 3864 6010 3888 6012
rect 3944 6010 3968 6012
rect 4024 6010 4048 6012
rect 4104 6010 4110 6012
rect 3864 5958 3866 6010
rect 4046 5958 4048 6010
rect 3802 5956 3808 5958
rect 3864 5956 3888 5958
rect 3944 5956 3968 5958
rect 4024 5956 4048 5958
rect 4104 5956 4110 5958
rect 3802 5947 4110 5956
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 1249 5468 1557 5477
rect 1249 5466 1255 5468
rect 1311 5466 1335 5468
rect 1391 5466 1415 5468
rect 1471 5466 1495 5468
rect 1551 5466 1557 5468
rect 1311 5414 1313 5466
rect 1493 5414 1495 5466
rect 1249 5412 1255 5414
rect 1311 5412 1335 5414
rect 1391 5412 1415 5414
rect 1471 5412 1495 5414
rect 1551 5412 1557 5414
rect 1249 5403 1557 5412
rect 2951 5468 3259 5477
rect 2951 5466 2957 5468
rect 3013 5466 3037 5468
rect 3093 5466 3117 5468
rect 3173 5466 3197 5468
rect 3253 5466 3259 5468
rect 3013 5414 3015 5466
rect 3195 5414 3197 5466
rect 2951 5412 2957 5414
rect 3013 5412 3037 5414
rect 3093 5412 3117 5414
rect 3173 5412 3197 5414
rect 3253 5412 3259 5414
rect 2951 5403 3259 5412
rect 3712 5370 3740 5714
rect 4172 5370 4200 6054
rect 4356 5846 4384 6054
rect 5000 5914 5028 7670
rect 6826 7600 6882 8000
rect 5504 7100 5812 7109
rect 5504 7098 5510 7100
rect 5566 7098 5590 7100
rect 5646 7098 5670 7100
rect 5726 7098 5750 7100
rect 5806 7098 5812 7100
rect 5566 7046 5568 7098
rect 5748 7046 5750 7098
rect 5504 7044 5510 7046
rect 5566 7044 5590 7046
rect 5646 7044 5670 7046
rect 5726 7044 5750 7046
rect 5806 7044 5812 7046
rect 5504 7035 5812 7044
rect 6840 7002 6868 7600
rect 7206 7100 7514 7109
rect 7206 7098 7212 7100
rect 7268 7098 7292 7100
rect 7348 7098 7372 7100
rect 7428 7098 7452 7100
rect 7508 7098 7514 7100
rect 7268 7046 7270 7098
rect 7450 7046 7452 7098
rect 7206 7044 7212 7046
rect 7268 7044 7292 7046
rect 7348 7044 7372 7046
rect 7428 7044 7452 7046
rect 7508 7044 7514 7046
rect 7206 7035 7514 7044
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 5276 5710 5304 6190
rect 5368 5846 5396 6598
rect 6355 6556 6663 6565
rect 6355 6554 6361 6556
rect 6417 6554 6441 6556
rect 6497 6554 6521 6556
rect 6577 6554 6601 6556
rect 6657 6554 6663 6556
rect 6417 6502 6419 6554
rect 6599 6502 6601 6554
rect 6355 6500 6361 6502
rect 6417 6500 6441 6502
rect 6497 6500 6521 6502
rect 6577 6500 6601 6502
rect 6657 6500 6663 6502
rect 6355 6491 6663 6500
rect 5504 6012 5812 6021
rect 5504 6010 5510 6012
rect 5566 6010 5590 6012
rect 5646 6010 5670 6012
rect 5726 6010 5750 6012
rect 5806 6010 5812 6012
rect 5566 5958 5568 6010
rect 5748 5958 5750 6010
rect 5504 5956 5510 5958
rect 5566 5956 5590 5958
rect 5646 5956 5670 5958
rect 5726 5956 5750 5958
rect 5806 5956 5812 5958
rect 5504 5947 5812 5956
rect 7206 6012 7514 6021
rect 7206 6010 7212 6012
rect 7268 6010 7292 6012
rect 7348 6010 7372 6012
rect 7428 6010 7452 6012
rect 7508 6010 7514 6012
rect 7268 5958 7270 6010
rect 7450 5958 7452 6010
rect 7206 5956 7212 5958
rect 7268 5956 7292 5958
rect 7348 5956 7372 5958
rect 7428 5956 7452 5958
rect 7508 5956 7514 5958
rect 7206 5947 7514 5956
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4653 5468 4961 5477
rect 4653 5466 4659 5468
rect 4715 5466 4739 5468
rect 4795 5466 4819 5468
rect 4875 5466 4899 5468
rect 4955 5466 4961 5468
rect 4715 5414 4717 5466
rect 4897 5414 4899 5466
rect 4653 5412 4659 5414
rect 4715 5412 4739 5414
rect 4795 5412 4819 5414
rect 4875 5412 4899 5414
rect 4955 5412 4961 5414
rect 4653 5403 4961 5412
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 5368 5030 5396 5782
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5234 5488 5646
rect 6355 5468 6663 5477
rect 6355 5466 6361 5468
rect 6417 5466 6441 5468
rect 6497 5466 6521 5468
rect 6577 5466 6601 5468
rect 6657 5466 6663 5468
rect 6417 5414 6419 5466
rect 6599 5414 6601 5466
rect 6355 5412 6361 5414
rect 6417 5412 6441 5414
rect 6497 5412 6521 5414
rect 6577 5412 6601 5414
rect 6657 5412 6663 5414
rect 6355 5403 6663 5412
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 2100 4924 2408 4933
rect 2100 4922 2106 4924
rect 2162 4922 2186 4924
rect 2242 4922 2266 4924
rect 2322 4922 2346 4924
rect 2402 4922 2408 4924
rect 2162 4870 2164 4922
rect 2344 4870 2346 4922
rect 2100 4868 2106 4870
rect 2162 4868 2186 4870
rect 2242 4868 2266 4870
rect 2322 4868 2346 4870
rect 2402 4868 2408 4870
rect 2100 4859 2408 4868
rect 3802 4924 4110 4933
rect 3802 4922 3808 4924
rect 3864 4922 3888 4924
rect 3944 4922 3968 4924
rect 4024 4922 4048 4924
rect 4104 4922 4110 4924
rect 3864 4870 3866 4922
rect 4046 4870 4048 4922
rect 3802 4868 3808 4870
rect 3864 4868 3888 4870
rect 3944 4868 3968 4870
rect 4024 4868 4048 4870
rect 4104 4868 4110 4870
rect 3802 4859 4110 4868
rect 5504 4924 5812 4933
rect 5504 4922 5510 4924
rect 5566 4922 5590 4924
rect 5646 4922 5670 4924
rect 5726 4922 5750 4924
rect 5806 4922 5812 4924
rect 5566 4870 5568 4922
rect 5748 4870 5750 4922
rect 5504 4868 5510 4870
rect 5566 4868 5590 4870
rect 5646 4868 5670 4870
rect 5726 4868 5750 4870
rect 5806 4868 5812 4870
rect 5504 4859 5812 4868
rect 7206 4924 7514 4933
rect 7206 4922 7212 4924
rect 7268 4922 7292 4924
rect 7348 4922 7372 4924
rect 7428 4922 7452 4924
rect 7508 4922 7514 4924
rect 7268 4870 7270 4922
rect 7450 4870 7452 4922
rect 7206 4868 7212 4870
rect 7268 4868 7292 4870
rect 7348 4868 7372 4870
rect 7428 4868 7452 4870
rect 7508 4868 7514 4870
rect 7206 4859 7514 4868
rect 1249 4380 1557 4389
rect 1249 4378 1255 4380
rect 1311 4378 1335 4380
rect 1391 4378 1415 4380
rect 1471 4378 1495 4380
rect 1551 4378 1557 4380
rect 1311 4326 1313 4378
rect 1493 4326 1495 4378
rect 1249 4324 1255 4326
rect 1311 4324 1335 4326
rect 1391 4324 1415 4326
rect 1471 4324 1495 4326
rect 1551 4324 1557 4326
rect 1249 4315 1557 4324
rect 2951 4380 3259 4389
rect 2951 4378 2957 4380
rect 3013 4378 3037 4380
rect 3093 4378 3117 4380
rect 3173 4378 3197 4380
rect 3253 4378 3259 4380
rect 3013 4326 3015 4378
rect 3195 4326 3197 4378
rect 2951 4324 2957 4326
rect 3013 4324 3037 4326
rect 3093 4324 3117 4326
rect 3173 4324 3197 4326
rect 3253 4324 3259 4326
rect 2951 4315 3259 4324
rect 4653 4380 4961 4389
rect 4653 4378 4659 4380
rect 4715 4378 4739 4380
rect 4795 4378 4819 4380
rect 4875 4378 4899 4380
rect 4955 4378 4961 4380
rect 4715 4326 4717 4378
rect 4897 4326 4899 4378
rect 4653 4324 4659 4326
rect 4715 4324 4739 4326
rect 4795 4324 4819 4326
rect 4875 4324 4899 4326
rect 4955 4324 4961 4326
rect 4653 4315 4961 4324
rect 6355 4380 6663 4389
rect 6355 4378 6361 4380
rect 6417 4378 6441 4380
rect 6497 4378 6521 4380
rect 6577 4378 6601 4380
rect 6657 4378 6663 4380
rect 6417 4326 6419 4378
rect 6599 4326 6601 4378
rect 6355 4324 6361 4326
rect 6417 4324 6441 4326
rect 6497 4324 6521 4326
rect 6577 4324 6601 4326
rect 6657 4324 6663 4326
rect 6355 4315 6663 4324
rect 2100 3836 2408 3845
rect 2100 3834 2106 3836
rect 2162 3834 2186 3836
rect 2242 3834 2266 3836
rect 2322 3834 2346 3836
rect 2402 3834 2408 3836
rect 2162 3782 2164 3834
rect 2344 3782 2346 3834
rect 2100 3780 2106 3782
rect 2162 3780 2186 3782
rect 2242 3780 2266 3782
rect 2322 3780 2346 3782
rect 2402 3780 2408 3782
rect 2100 3771 2408 3780
rect 3802 3836 4110 3845
rect 3802 3834 3808 3836
rect 3864 3834 3888 3836
rect 3944 3834 3968 3836
rect 4024 3834 4048 3836
rect 4104 3834 4110 3836
rect 3864 3782 3866 3834
rect 4046 3782 4048 3834
rect 3802 3780 3808 3782
rect 3864 3780 3888 3782
rect 3944 3780 3968 3782
rect 4024 3780 4048 3782
rect 4104 3780 4110 3782
rect 3802 3771 4110 3780
rect 5504 3836 5812 3845
rect 5504 3834 5510 3836
rect 5566 3834 5590 3836
rect 5646 3834 5670 3836
rect 5726 3834 5750 3836
rect 5806 3834 5812 3836
rect 5566 3782 5568 3834
rect 5748 3782 5750 3834
rect 5504 3780 5510 3782
rect 5566 3780 5590 3782
rect 5646 3780 5670 3782
rect 5726 3780 5750 3782
rect 5806 3780 5812 3782
rect 5504 3771 5812 3780
rect 7206 3836 7514 3845
rect 7206 3834 7212 3836
rect 7268 3834 7292 3836
rect 7348 3834 7372 3836
rect 7428 3834 7452 3836
rect 7508 3834 7514 3836
rect 7268 3782 7270 3834
rect 7450 3782 7452 3834
rect 7206 3780 7212 3782
rect 7268 3780 7292 3782
rect 7348 3780 7372 3782
rect 7428 3780 7452 3782
rect 7508 3780 7514 3782
rect 7206 3771 7514 3780
rect 1249 3292 1557 3301
rect 1249 3290 1255 3292
rect 1311 3290 1335 3292
rect 1391 3290 1415 3292
rect 1471 3290 1495 3292
rect 1551 3290 1557 3292
rect 1311 3238 1313 3290
rect 1493 3238 1495 3290
rect 1249 3236 1255 3238
rect 1311 3236 1335 3238
rect 1391 3236 1415 3238
rect 1471 3236 1495 3238
rect 1551 3236 1557 3238
rect 1249 3227 1557 3236
rect 2951 3292 3259 3301
rect 2951 3290 2957 3292
rect 3013 3290 3037 3292
rect 3093 3290 3117 3292
rect 3173 3290 3197 3292
rect 3253 3290 3259 3292
rect 3013 3238 3015 3290
rect 3195 3238 3197 3290
rect 2951 3236 2957 3238
rect 3013 3236 3037 3238
rect 3093 3236 3117 3238
rect 3173 3236 3197 3238
rect 3253 3236 3259 3238
rect 2951 3227 3259 3236
rect 4653 3292 4961 3301
rect 4653 3290 4659 3292
rect 4715 3290 4739 3292
rect 4795 3290 4819 3292
rect 4875 3290 4899 3292
rect 4955 3290 4961 3292
rect 4715 3238 4717 3290
rect 4897 3238 4899 3290
rect 4653 3236 4659 3238
rect 4715 3236 4739 3238
rect 4795 3236 4819 3238
rect 4875 3236 4899 3238
rect 4955 3236 4961 3238
rect 4653 3227 4961 3236
rect 6355 3292 6663 3301
rect 6355 3290 6361 3292
rect 6417 3290 6441 3292
rect 6497 3290 6521 3292
rect 6577 3290 6601 3292
rect 6657 3290 6663 3292
rect 6417 3238 6419 3290
rect 6599 3238 6601 3290
rect 6355 3236 6361 3238
rect 6417 3236 6441 3238
rect 6497 3236 6521 3238
rect 6577 3236 6601 3238
rect 6657 3236 6663 3238
rect 6355 3227 6663 3236
rect 2100 2748 2408 2757
rect 2100 2746 2106 2748
rect 2162 2746 2186 2748
rect 2242 2746 2266 2748
rect 2322 2746 2346 2748
rect 2402 2746 2408 2748
rect 2162 2694 2164 2746
rect 2344 2694 2346 2746
rect 2100 2692 2106 2694
rect 2162 2692 2186 2694
rect 2242 2692 2266 2694
rect 2322 2692 2346 2694
rect 2402 2692 2408 2694
rect 2100 2683 2408 2692
rect 3802 2748 4110 2757
rect 3802 2746 3808 2748
rect 3864 2746 3888 2748
rect 3944 2746 3968 2748
rect 4024 2746 4048 2748
rect 4104 2746 4110 2748
rect 3864 2694 3866 2746
rect 4046 2694 4048 2746
rect 3802 2692 3808 2694
rect 3864 2692 3888 2694
rect 3944 2692 3968 2694
rect 4024 2692 4048 2694
rect 4104 2692 4110 2694
rect 3802 2683 4110 2692
rect 5504 2748 5812 2757
rect 5504 2746 5510 2748
rect 5566 2746 5590 2748
rect 5646 2746 5670 2748
rect 5726 2746 5750 2748
rect 5806 2746 5812 2748
rect 5566 2694 5568 2746
rect 5748 2694 5750 2746
rect 5504 2692 5510 2694
rect 5566 2692 5590 2694
rect 5646 2692 5670 2694
rect 5726 2692 5750 2694
rect 5806 2692 5812 2694
rect 5504 2683 5812 2692
rect 7206 2748 7514 2757
rect 7206 2746 7212 2748
rect 7268 2746 7292 2748
rect 7348 2746 7372 2748
rect 7428 2746 7452 2748
rect 7508 2746 7514 2748
rect 7268 2694 7270 2746
rect 7450 2694 7452 2746
rect 7206 2692 7212 2694
rect 7268 2692 7292 2694
rect 7348 2692 7372 2694
rect 7428 2692 7452 2694
rect 7508 2692 7514 2694
rect 7206 2683 7514 2692
rect 1249 2204 1557 2213
rect 1249 2202 1255 2204
rect 1311 2202 1335 2204
rect 1391 2202 1415 2204
rect 1471 2202 1495 2204
rect 1551 2202 1557 2204
rect 1311 2150 1313 2202
rect 1493 2150 1495 2202
rect 1249 2148 1255 2150
rect 1311 2148 1335 2150
rect 1391 2148 1415 2150
rect 1471 2148 1495 2150
rect 1551 2148 1557 2150
rect 1249 2139 1557 2148
rect 2951 2204 3259 2213
rect 2951 2202 2957 2204
rect 3013 2202 3037 2204
rect 3093 2202 3117 2204
rect 3173 2202 3197 2204
rect 3253 2202 3259 2204
rect 3013 2150 3015 2202
rect 3195 2150 3197 2202
rect 2951 2148 2957 2150
rect 3013 2148 3037 2150
rect 3093 2148 3117 2150
rect 3173 2148 3197 2150
rect 3253 2148 3259 2150
rect 2951 2139 3259 2148
rect 4653 2204 4961 2213
rect 4653 2202 4659 2204
rect 4715 2202 4739 2204
rect 4795 2202 4819 2204
rect 4875 2202 4899 2204
rect 4955 2202 4961 2204
rect 4715 2150 4717 2202
rect 4897 2150 4899 2202
rect 4653 2148 4659 2150
rect 4715 2148 4739 2150
rect 4795 2148 4819 2150
rect 4875 2148 4899 2150
rect 4955 2148 4961 2150
rect 4653 2139 4961 2148
rect 6355 2204 6663 2213
rect 6355 2202 6361 2204
rect 6417 2202 6441 2204
rect 6497 2202 6521 2204
rect 6577 2202 6601 2204
rect 6657 2202 6663 2204
rect 6417 2150 6419 2202
rect 6599 2150 6601 2202
rect 6355 2148 6361 2150
rect 6417 2148 6441 2150
rect 6497 2148 6521 2150
rect 6577 2148 6601 2150
rect 6657 2148 6663 2150
rect 6355 2139 6663 2148
rect 2100 1660 2408 1669
rect 2100 1658 2106 1660
rect 2162 1658 2186 1660
rect 2242 1658 2266 1660
rect 2322 1658 2346 1660
rect 2402 1658 2408 1660
rect 2162 1606 2164 1658
rect 2344 1606 2346 1658
rect 2100 1604 2106 1606
rect 2162 1604 2186 1606
rect 2242 1604 2266 1606
rect 2322 1604 2346 1606
rect 2402 1604 2408 1606
rect 2100 1595 2408 1604
rect 3802 1660 4110 1669
rect 3802 1658 3808 1660
rect 3864 1658 3888 1660
rect 3944 1658 3968 1660
rect 4024 1658 4048 1660
rect 4104 1658 4110 1660
rect 3864 1606 3866 1658
rect 4046 1606 4048 1658
rect 3802 1604 3808 1606
rect 3864 1604 3888 1606
rect 3944 1604 3968 1606
rect 4024 1604 4048 1606
rect 4104 1604 4110 1606
rect 3802 1595 4110 1604
rect 5504 1660 5812 1669
rect 5504 1658 5510 1660
rect 5566 1658 5590 1660
rect 5646 1658 5670 1660
rect 5726 1658 5750 1660
rect 5806 1658 5812 1660
rect 5566 1606 5568 1658
rect 5748 1606 5750 1658
rect 5504 1604 5510 1606
rect 5566 1604 5590 1606
rect 5646 1604 5670 1606
rect 5726 1604 5750 1606
rect 5806 1604 5812 1606
rect 5504 1595 5812 1604
rect 7206 1660 7514 1669
rect 7206 1658 7212 1660
rect 7268 1658 7292 1660
rect 7348 1658 7372 1660
rect 7428 1658 7452 1660
rect 7508 1658 7514 1660
rect 7268 1606 7270 1658
rect 7450 1606 7452 1658
rect 7206 1604 7212 1606
rect 7268 1604 7292 1606
rect 7348 1604 7372 1606
rect 7428 1604 7452 1606
rect 7508 1604 7514 1606
rect 7206 1595 7514 1604
rect 1249 1116 1557 1125
rect 1249 1114 1255 1116
rect 1311 1114 1335 1116
rect 1391 1114 1415 1116
rect 1471 1114 1495 1116
rect 1551 1114 1557 1116
rect 1311 1062 1313 1114
rect 1493 1062 1495 1114
rect 1249 1060 1255 1062
rect 1311 1060 1335 1062
rect 1391 1060 1415 1062
rect 1471 1060 1495 1062
rect 1551 1060 1557 1062
rect 1249 1051 1557 1060
rect 2951 1116 3259 1125
rect 2951 1114 2957 1116
rect 3013 1114 3037 1116
rect 3093 1114 3117 1116
rect 3173 1114 3197 1116
rect 3253 1114 3259 1116
rect 3013 1062 3015 1114
rect 3195 1062 3197 1114
rect 2951 1060 2957 1062
rect 3013 1060 3037 1062
rect 3093 1060 3117 1062
rect 3173 1060 3197 1062
rect 3253 1060 3259 1062
rect 2951 1051 3259 1060
rect 4653 1116 4961 1125
rect 4653 1114 4659 1116
rect 4715 1114 4739 1116
rect 4795 1114 4819 1116
rect 4875 1114 4899 1116
rect 4955 1114 4961 1116
rect 4715 1062 4717 1114
rect 4897 1062 4899 1114
rect 4653 1060 4659 1062
rect 4715 1060 4739 1062
rect 4795 1060 4819 1062
rect 4875 1060 4899 1062
rect 4955 1060 4961 1062
rect 4653 1051 4961 1060
rect 6355 1116 6663 1125
rect 6355 1114 6361 1116
rect 6417 1114 6441 1116
rect 6497 1114 6521 1116
rect 6577 1114 6601 1116
rect 6657 1114 6663 1116
rect 6417 1062 6419 1114
rect 6599 1062 6601 1114
rect 6355 1060 6361 1062
rect 6417 1060 6441 1062
rect 6497 1060 6521 1062
rect 6577 1060 6601 1062
rect 6657 1060 6663 1062
rect 6355 1051 6663 1060
rect 2100 572 2408 581
rect 2100 570 2106 572
rect 2162 570 2186 572
rect 2242 570 2266 572
rect 2322 570 2346 572
rect 2402 570 2408 572
rect 2162 518 2164 570
rect 2344 518 2346 570
rect 2100 516 2106 518
rect 2162 516 2186 518
rect 2242 516 2266 518
rect 2322 516 2346 518
rect 2402 516 2408 518
rect 2100 507 2408 516
rect 3802 572 4110 581
rect 3802 570 3808 572
rect 3864 570 3888 572
rect 3944 570 3968 572
rect 4024 570 4048 572
rect 4104 570 4110 572
rect 3864 518 3866 570
rect 4046 518 4048 570
rect 3802 516 3808 518
rect 3864 516 3888 518
rect 3944 516 3968 518
rect 4024 516 4048 518
rect 4104 516 4110 518
rect 3802 507 4110 516
rect 5504 572 5812 581
rect 5504 570 5510 572
rect 5566 570 5590 572
rect 5646 570 5670 572
rect 5726 570 5750 572
rect 5806 570 5812 572
rect 5566 518 5568 570
rect 5748 518 5750 570
rect 5504 516 5510 518
rect 5566 516 5590 518
rect 5646 516 5670 518
rect 5726 516 5750 518
rect 5806 516 5812 518
rect 5504 507 5812 516
rect 7206 572 7514 581
rect 7206 570 7212 572
rect 7268 570 7292 572
rect 7348 570 7372 572
rect 7428 570 7452 572
rect 7508 570 7514 572
rect 7268 518 7270 570
rect 7450 518 7452 570
rect 7206 516 7212 518
rect 7268 516 7292 518
rect 7348 516 7372 518
rect 7428 516 7452 518
rect 7508 516 7514 518
rect 7206 507 7514 516
<< via2 >>
rect 1255 6554 1311 6556
rect 1335 6554 1391 6556
rect 1415 6554 1471 6556
rect 1495 6554 1551 6556
rect 1255 6502 1301 6554
rect 1301 6502 1311 6554
rect 1335 6502 1365 6554
rect 1365 6502 1377 6554
rect 1377 6502 1391 6554
rect 1415 6502 1429 6554
rect 1429 6502 1441 6554
rect 1441 6502 1471 6554
rect 1495 6502 1505 6554
rect 1505 6502 1551 6554
rect 1255 6500 1311 6502
rect 1335 6500 1391 6502
rect 1415 6500 1471 6502
rect 1495 6500 1551 6502
rect 2106 7098 2162 7100
rect 2186 7098 2242 7100
rect 2266 7098 2322 7100
rect 2346 7098 2402 7100
rect 2106 7046 2152 7098
rect 2152 7046 2162 7098
rect 2186 7046 2216 7098
rect 2216 7046 2228 7098
rect 2228 7046 2242 7098
rect 2266 7046 2280 7098
rect 2280 7046 2292 7098
rect 2292 7046 2322 7098
rect 2346 7046 2356 7098
rect 2356 7046 2402 7098
rect 2106 7044 2162 7046
rect 2186 7044 2242 7046
rect 2266 7044 2322 7046
rect 2346 7044 2402 7046
rect 3808 7098 3864 7100
rect 3888 7098 3944 7100
rect 3968 7098 4024 7100
rect 4048 7098 4104 7100
rect 3808 7046 3854 7098
rect 3854 7046 3864 7098
rect 3888 7046 3918 7098
rect 3918 7046 3930 7098
rect 3930 7046 3944 7098
rect 3968 7046 3982 7098
rect 3982 7046 3994 7098
rect 3994 7046 4024 7098
rect 4048 7046 4058 7098
rect 4058 7046 4104 7098
rect 3808 7044 3864 7046
rect 3888 7044 3944 7046
rect 3968 7044 4024 7046
rect 4048 7044 4104 7046
rect 2957 6554 3013 6556
rect 3037 6554 3093 6556
rect 3117 6554 3173 6556
rect 3197 6554 3253 6556
rect 2957 6502 3003 6554
rect 3003 6502 3013 6554
rect 3037 6502 3067 6554
rect 3067 6502 3079 6554
rect 3079 6502 3093 6554
rect 3117 6502 3131 6554
rect 3131 6502 3143 6554
rect 3143 6502 3173 6554
rect 3197 6502 3207 6554
rect 3207 6502 3253 6554
rect 2957 6500 3013 6502
rect 3037 6500 3093 6502
rect 3117 6500 3173 6502
rect 3197 6500 3253 6502
rect 4659 6554 4715 6556
rect 4739 6554 4795 6556
rect 4819 6554 4875 6556
rect 4899 6554 4955 6556
rect 4659 6502 4705 6554
rect 4705 6502 4715 6554
rect 4739 6502 4769 6554
rect 4769 6502 4781 6554
rect 4781 6502 4795 6554
rect 4819 6502 4833 6554
rect 4833 6502 4845 6554
rect 4845 6502 4875 6554
rect 4899 6502 4909 6554
rect 4909 6502 4955 6554
rect 4659 6500 4715 6502
rect 4739 6500 4795 6502
rect 4819 6500 4875 6502
rect 4899 6500 4955 6502
rect 2106 6010 2162 6012
rect 2186 6010 2242 6012
rect 2266 6010 2322 6012
rect 2346 6010 2402 6012
rect 2106 5958 2152 6010
rect 2152 5958 2162 6010
rect 2186 5958 2216 6010
rect 2216 5958 2228 6010
rect 2228 5958 2242 6010
rect 2266 5958 2280 6010
rect 2280 5958 2292 6010
rect 2292 5958 2322 6010
rect 2346 5958 2356 6010
rect 2356 5958 2402 6010
rect 2106 5956 2162 5958
rect 2186 5956 2242 5958
rect 2266 5956 2322 5958
rect 2346 5956 2402 5958
rect 3808 6010 3864 6012
rect 3888 6010 3944 6012
rect 3968 6010 4024 6012
rect 4048 6010 4104 6012
rect 3808 5958 3854 6010
rect 3854 5958 3864 6010
rect 3888 5958 3918 6010
rect 3918 5958 3930 6010
rect 3930 5958 3944 6010
rect 3968 5958 3982 6010
rect 3982 5958 3994 6010
rect 3994 5958 4024 6010
rect 4048 5958 4058 6010
rect 4058 5958 4104 6010
rect 3808 5956 3864 5958
rect 3888 5956 3944 5958
rect 3968 5956 4024 5958
rect 4048 5956 4104 5958
rect 1255 5466 1311 5468
rect 1335 5466 1391 5468
rect 1415 5466 1471 5468
rect 1495 5466 1551 5468
rect 1255 5414 1301 5466
rect 1301 5414 1311 5466
rect 1335 5414 1365 5466
rect 1365 5414 1377 5466
rect 1377 5414 1391 5466
rect 1415 5414 1429 5466
rect 1429 5414 1441 5466
rect 1441 5414 1471 5466
rect 1495 5414 1505 5466
rect 1505 5414 1551 5466
rect 1255 5412 1311 5414
rect 1335 5412 1391 5414
rect 1415 5412 1471 5414
rect 1495 5412 1551 5414
rect 2957 5466 3013 5468
rect 3037 5466 3093 5468
rect 3117 5466 3173 5468
rect 3197 5466 3253 5468
rect 2957 5414 3003 5466
rect 3003 5414 3013 5466
rect 3037 5414 3067 5466
rect 3067 5414 3079 5466
rect 3079 5414 3093 5466
rect 3117 5414 3131 5466
rect 3131 5414 3143 5466
rect 3143 5414 3173 5466
rect 3197 5414 3207 5466
rect 3207 5414 3253 5466
rect 2957 5412 3013 5414
rect 3037 5412 3093 5414
rect 3117 5412 3173 5414
rect 3197 5412 3253 5414
rect 5510 7098 5566 7100
rect 5590 7098 5646 7100
rect 5670 7098 5726 7100
rect 5750 7098 5806 7100
rect 5510 7046 5556 7098
rect 5556 7046 5566 7098
rect 5590 7046 5620 7098
rect 5620 7046 5632 7098
rect 5632 7046 5646 7098
rect 5670 7046 5684 7098
rect 5684 7046 5696 7098
rect 5696 7046 5726 7098
rect 5750 7046 5760 7098
rect 5760 7046 5806 7098
rect 5510 7044 5566 7046
rect 5590 7044 5646 7046
rect 5670 7044 5726 7046
rect 5750 7044 5806 7046
rect 7212 7098 7268 7100
rect 7292 7098 7348 7100
rect 7372 7098 7428 7100
rect 7452 7098 7508 7100
rect 7212 7046 7258 7098
rect 7258 7046 7268 7098
rect 7292 7046 7322 7098
rect 7322 7046 7334 7098
rect 7334 7046 7348 7098
rect 7372 7046 7386 7098
rect 7386 7046 7398 7098
rect 7398 7046 7428 7098
rect 7452 7046 7462 7098
rect 7462 7046 7508 7098
rect 7212 7044 7268 7046
rect 7292 7044 7348 7046
rect 7372 7044 7428 7046
rect 7452 7044 7508 7046
rect 6361 6554 6417 6556
rect 6441 6554 6497 6556
rect 6521 6554 6577 6556
rect 6601 6554 6657 6556
rect 6361 6502 6407 6554
rect 6407 6502 6417 6554
rect 6441 6502 6471 6554
rect 6471 6502 6483 6554
rect 6483 6502 6497 6554
rect 6521 6502 6535 6554
rect 6535 6502 6547 6554
rect 6547 6502 6577 6554
rect 6601 6502 6611 6554
rect 6611 6502 6657 6554
rect 6361 6500 6417 6502
rect 6441 6500 6497 6502
rect 6521 6500 6577 6502
rect 6601 6500 6657 6502
rect 5510 6010 5566 6012
rect 5590 6010 5646 6012
rect 5670 6010 5726 6012
rect 5750 6010 5806 6012
rect 5510 5958 5556 6010
rect 5556 5958 5566 6010
rect 5590 5958 5620 6010
rect 5620 5958 5632 6010
rect 5632 5958 5646 6010
rect 5670 5958 5684 6010
rect 5684 5958 5696 6010
rect 5696 5958 5726 6010
rect 5750 5958 5760 6010
rect 5760 5958 5806 6010
rect 5510 5956 5566 5958
rect 5590 5956 5646 5958
rect 5670 5956 5726 5958
rect 5750 5956 5806 5958
rect 7212 6010 7268 6012
rect 7292 6010 7348 6012
rect 7372 6010 7428 6012
rect 7452 6010 7508 6012
rect 7212 5958 7258 6010
rect 7258 5958 7268 6010
rect 7292 5958 7322 6010
rect 7322 5958 7334 6010
rect 7334 5958 7348 6010
rect 7372 5958 7386 6010
rect 7386 5958 7398 6010
rect 7398 5958 7428 6010
rect 7452 5958 7462 6010
rect 7462 5958 7508 6010
rect 7212 5956 7268 5958
rect 7292 5956 7348 5958
rect 7372 5956 7428 5958
rect 7452 5956 7508 5958
rect 4659 5466 4715 5468
rect 4739 5466 4795 5468
rect 4819 5466 4875 5468
rect 4899 5466 4955 5468
rect 4659 5414 4705 5466
rect 4705 5414 4715 5466
rect 4739 5414 4769 5466
rect 4769 5414 4781 5466
rect 4781 5414 4795 5466
rect 4819 5414 4833 5466
rect 4833 5414 4845 5466
rect 4845 5414 4875 5466
rect 4899 5414 4909 5466
rect 4909 5414 4955 5466
rect 4659 5412 4715 5414
rect 4739 5412 4795 5414
rect 4819 5412 4875 5414
rect 4899 5412 4955 5414
rect 6361 5466 6417 5468
rect 6441 5466 6497 5468
rect 6521 5466 6577 5468
rect 6601 5466 6657 5468
rect 6361 5414 6407 5466
rect 6407 5414 6417 5466
rect 6441 5414 6471 5466
rect 6471 5414 6483 5466
rect 6483 5414 6497 5466
rect 6521 5414 6535 5466
rect 6535 5414 6547 5466
rect 6547 5414 6577 5466
rect 6601 5414 6611 5466
rect 6611 5414 6657 5466
rect 6361 5412 6417 5414
rect 6441 5412 6497 5414
rect 6521 5412 6577 5414
rect 6601 5412 6657 5414
rect 2106 4922 2162 4924
rect 2186 4922 2242 4924
rect 2266 4922 2322 4924
rect 2346 4922 2402 4924
rect 2106 4870 2152 4922
rect 2152 4870 2162 4922
rect 2186 4870 2216 4922
rect 2216 4870 2228 4922
rect 2228 4870 2242 4922
rect 2266 4870 2280 4922
rect 2280 4870 2292 4922
rect 2292 4870 2322 4922
rect 2346 4870 2356 4922
rect 2356 4870 2402 4922
rect 2106 4868 2162 4870
rect 2186 4868 2242 4870
rect 2266 4868 2322 4870
rect 2346 4868 2402 4870
rect 3808 4922 3864 4924
rect 3888 4922 3944 4924
rect 3968 4922 4024 4924
rect 4048 4922 4104 4924
rect 3808 4870 3854 4922
rect 3854 4870 3864 4922
rect 3888 4870 3918 4922
rect 3918 4870 3930 4922
rect 3930 4870 3944 4922
rect 3968 4870 3982 4922
rect 3982 4870 3994 4922
rect 3994 4870 4024 4922
rect 4048 4870 4058 4922
rect 4058 4870 4104 4922
rect 3808 4868 3864 4870
rect 3888 4868 3944 4870
rect 3968 4868 4024 4870
rect 4048 4868 4104 4870
rect 5510 4922 5566 4924
rect 5590 4922 5646 4924
rect 5670 4922 5726 4924
rect 5750 4922 5806 4924
rect 5510 4870 5556 4922
rect 5556 4870 5566 4922
rect 5590 4870 5620 4922
rect 5620 4870 5632 4922
rect 5632 4870 5646 4922
rect 5670 4870 5684 4922
rect 5684 4870 5696 4922
rect 5696 4870 5726 4922
rect 5750 4870 5760 4922
rect 5760 4870 5806 4922
rect 5510 4868 5566 4870
rect 5590 4868 5646 4870
rect 5670 4868 5726 4870
rect 5750 4868 5806 4870
rect 7212 4922 7268 4924
rect 7292 4922 7348 4924
rect 7372 4922 7428 4924
rect 7452 4922 7508 4924
rect 7212 4870 7258 4922
rect 7258 4870 7268 4922
rect 7292 4870 7322 4922
rect 7322 4870 7334 4922
rect 7334 4870 7348 4922
rect 7372 4870 7386 4922
rect 7386 4870 7398 4922
rect 7398 4870 7428 4922
rect 7452 4870 7462 4922
rect 7462 4870 7508 4922
rect 7212 4868 7268 4870
rect 7292 4868 7348 4870
rect 7372 4868 7428 4870
rect 7452 4868 7508 4870
rect 1255 4378 1311 4380
rect 1335 4378 1391 4380
rect 1415 4378 1471 4380
rect 1495 4378 1551 4380
rect 1255 4326 1301 4378
rect 1301 4326 1311 4378
rect 1335 4326 1365 4378
rect 1365 4326 1377 4378
rect 1377 4326 1391 4378
rect 1415 4326 1429 4378
rect 1429 4326 1441 4378
rect 1441 4326 1471 4378
rect 1495 4326 1505 4378
rect 1505 4326 1551 4378
rect 1255 4324 1311 4326
rect 1335 4324 1391 4326
rect 1415 4324 1471 4326
rect 1495 4324 1551 4326
rect 2957 4378 3013 4380
rect 3037 4378 3093 4380
rect 3117 4378 3173 4380
rect 3197 4378 3253 4380
rect 2957 4326 3003 4378
rect 3003 4326 3013 4378
rect 3037 4326 3067 4378
rect 3067 4326 3079 4378
rect 3079 4326 3093 4378
rect 3117 4326 3131 4378
rect 3131 4326 3143 4378
rect 3143 4326 3173 4378
rect 3197 4326 3207 4378
rect 3207 4326 3253 4378
rect 2957 4324 3013 4326
rect 3037 4324 3093 4326
rect 3117 4324 3173 4326
rect 3197 4324 3253 4326
rect 4659 4378 4715 4380
rect 4739 4378 4795 4380
rect 4819 4378 4875 4380
rect 4899 4378 4955 4380
rect 4659 4326 4705 4378
rect 4705 4326 4715 4378
rect 4739 4326 4769 4378
rect 4769 4326 4781 4378
rect 4781 4326 4795 4378
rect 4819 4326 4833 4378
rect 4833 4326 4845 4378
rect 4845 4326 4875 4378
rect 4899 4326 4909 4378
rect 4909 4326 4955 4378
rect 4659 4324 4715 4326
rect 4739 4324 4795 4326
rect 4819 4324 4875 4326
rect 4899 4324 4955 4326
rect 6361 4378 6417 4380
rect 6441 4378 6497 4380
rect 6521 4378 6577 4380
rect 6601 4378 6657 4380
rect 6361 4326 6407 4378
rect 6407 4326 6417 4378
rect 6441 4326 6471 4378
rect 6471 4326 6483 4378
rect 6483 4326 6497 4378
rect 6521 4326 6535 4378
rect 6535 4326 6547 4378
rect 6547 4326 6577 4378
rect 6601 4326 6611 4378
rect 6611 4326 6657 4378
rect 6361 4324 6417 4326
rect 6441 4324 6497 4326
rect 6521 4324 6577 4326
rect 6601 4324 6657 4326
rect 2106 3834 2162 3836
rect 2186 3834 2242 3836
rect 2266 3834 2322 3836
rect 2346 3834 2402 3836
rect 2106 3782 2152 3834
rect 2152 3782 2162 3834
rect 2186 3782 2216 3834
rect 2216 3782 2228 3834
rect 2228 3782 2242 3834
rect 2266 3782 2280 3834
rect 2280 3782 2292 3834
rect 2292 3782 2322 3834
rect 2346 3782 2356 3834
rect 2356 3782 2402 3834
rect 2106 3780 2162 3782
rect 2186 3780 2242 3782
rect 2266 3780 2322 3782
rect 2346 3780 2402 3782
rect 3808 3834 3864 3836
rect 3888 3834 3944 3836
rect 3968 3834 4024 3836
rect 4048 3834 4104 3836
rect 3808 3782 3854 3834
rect 3854 3782 3864 3834
rect 3888 3782 3918 3834
rect 3918 3782 3930 3834
rect 3930 3782 3944 3834
rect 3968 3782 3982 3834
rect 3982 3782 3994 3834
rect 3994 3782 4024 3834
rect 4048 3782 4058 3834
rect 4058 3782 4104 3834
rect 3808 3780 3864 3782
rect 3888 3780 3944 3782
rect 3968 3780 4024 3782
rect 4048 3780 4104 3782
rect 5510 3834 5566 3836
rect 5590 3834 5646 3836
rect 5670 3834 5726 3836
rect 5750 3834 5806 3836
rect 5510 3782 5556 3834
rect 5556 3782 5566 3834
rect 5590 3782 5620 3834
rect 5620 3782 5632 3834
rect 5632 3782 5646 3834
rect 5670 3782 5684 3834
rect 5684 3782 5696 3834
rect 5696 3782 5726 3834
rect 5750 3782 5760 3834
rect 5760 3782 5806 3834
rect 5510 3780 5566 3782
rect 5590 3780 5646 3782
rect 5670 3780 5726 3782
rect 5750 3780 5806 3782
rect 7212 3834 7268 3836
rect 7292 3834 7348 3836
rect 7372 3834 7428 3836
rect 7452 3834 7508 3836
rect 7212 3782 7258 3834
rect 7258 3782 7268 3834
rect 7292 3782 7322 3834
rect 7322 3782 7334 3834
rect 7334 3782 7348 3834
rect 7372 3782 7386 3834
rect 7386 3782 7398 3834
rect 7398 3782 7428 3834
rect 7452 3782 7462 3834
rect 7462 3782 7508 3834
rect 7212 3780 7268 3782
rect 7292 3780 7348 3782
rect 7372 3780 7428 3782
rect 7452 3780 7508 3782
rect 1255 3290 1311 3292
rect 1335 3290 1391 3292
rect 1415 3290 1471 3292
rect 1495 3290 1551 3292
rect 1255 3238 1301 3290
rect 1301 3238 1311 3290
rect 1335 3238 1365 3290
rect 1365 3238 1377 3290
rect 1377 3238 1391 3290
rect 1415 3238 1429 3290
rect 1429 3238 1441 3290
rect 1441 3238 1471 3290
rect 1495 3238 1505 3290
rect 1505 3238 1551 3290
rect 1255 3236 1311 3238
rect 1335 3236 1391 3238
rect 1415 3236 1471 3238
rect 1495 3236 1551 3238
rect 2957 3290 3013 3292
rect 3037 3290 3093 3292
rect 3117 3290 3173 3292
rect 3197 3290 3253 3292
rect 2957 3238 3003 3290
rect 3003 3238 3013 3290
rect 3037 3238 3067 3290
rect 3067 3238 3079 3290
rect 3079 3238 3093 3290
rect 3117 3238 3131 3290
rect 3131 3238 3143 3290
rect 3143 3238 3173 3290
rect 3197 3238 3207 3290
rect 3207 3238 3253 3290
rect 2957 3236 3013 3238
rect 3037 3236 3093 3238
rect 3117 3236 3173 3238
rect 3197 3236 3253 3238
rect 4659 3290 4715 3292
rect 4739 3290 4795 3292
rect 4819 3290 4875 3292
rect 4899 3290 4955 3292
rect 4659 3238 4705 3290
rect 4705 3238 4715 3290
rect 4739 3238 4769 3290
rect 4769 3238 4781 3290
rect 4781 3238 4795 3290
rect 4819 3238 4833 3290
rect 4833 3238 4845 3290
rect 4845 3238 4875 3290
rect 4899 3238 4909 3290
rect 4909 3238 4955 3290
rect 4659 3236 4715 3238
rect 4739 3236 4795 3238
rect 4819 3236 4875 3238
rect 4899 3236 4955 3238
rect 6361 3290 6417 3292
rect 6441 3290 6497 3292
rect 6521 3290 6577 3292
rect 6601 3290 6657 3292
rect 6361 3238 6407 3290
rect 6407 3238 6417 3290
rect 6441 3238 6471 3290
rect 6471 3238 6483 3290
rect 6483 3238 6497 3290
rect 6521 3238 6535 3290
rect 6535 3238 6547 3290
rect 6547 3238 6577 3290
rect 6601 3238 6611 3290
rect 6611 3238 6657 3290
rect 6361 3236 6417 3238
rect 6441 3236 6497 3238
rect 6521 3236 6577 3238
rect 6601 3236 6657 3238
rect 2106 2746 2162 2748
rect 2186 2746 2242 2748
rect 2266 2746 2322 2748
rect 2346 2746 2402 2748
rect 2106 2694 2152 2746
rect 2152 2694 2162 2746
rect 2186 2694 2216 2746
rect 2216 2694 2228 2746
rect 2228 2694 2242 2746
rect 2266 2694 2280 2746
rect 2280 2694 2292 2746
rect 2292 2694 2322 2746
rect 2346 2694 2356 2746
rect 2356 2694 2402 2746
rect 2106 2692 2162 2694
rect 2186 2692 2242 2694
rect 2266 2692 2322 2694
rect 2346 2692 2402 2694
rect 3808 2746 3864 2748
rect 3888 2746 3944 2748
rect 3968 2746 4024 2748
rect 4048 2746 4104 2748
rect 3808 2694 3854 2746
rect 3854 2694 3864 2746
rect 3888 2694 3918 2746
rect 3918 2694 3930 2746
rect 3930 2694 3944 2746
rect 3968 2694 3982 2746
rect 3982 2694 3994 2746
rect 3994 2694 4024 2746
rect 4048 2694 4058 2746
rect 4058 2694 4104 2746
rect 3808 2692 3864 2694
rect 3888 2692 3944 2694
rect 3968 2692 4024 2694
rect 4048 2692 4104 2694
rect 5510 2746 5566 2748
rect 5590 2746 5646 2748
rect 5670 2746 5726 2748
rect 5750 2746 5806 2748
rect 5510 2694 5556 2746
rect 5556 2694 5566 2746
rect 5590 2694 5620 2746
rect 5620 2694 5632 2746
rect 5632 2694 5646 2746
rect 5670 2694 5684 2746
rect 5684 2694 5696 2746
rect 5696 2694 5726 2746
rect 5750 2694 5760 2746
rect 5760 2694 5806 2746
rect 5510 2692 5566 2694
rect 5590 2692 5646 2694
rect 5670 2692 5726 2694
rect 5750 2692 5806 2694
rect 7212 2746 7268 2748
rect 7292 2746 7348 2748
rect 7372 2746 7428 2748
rect 7452 2746 7508 2748
rect 7212 2694 7258 2746
rect 7258 2694 7268 2746
rect 7292 2694 7322 2746
rect 7322 2694 7334 2746
rect 7334 2694 7348 2746
rect 7372 2694 7386 2746
rect 7386 2694 7398 2746
rect 7398 2694 7428 2746
rect 7452 2694 7462 2746
rect 7462 2694 7508 2746
rect 7212 2692 7268 2694
rect 7292 2692 7348 2694
rect 7372 2692 7428 2694
rect 7452 2692 7508 2694
rect 1255 2202 1311 2204
rect 1335 2202 1391 2204
rect 1415 2202 1471 2204
rect 1495 2202 1551 2204
rect 1255 2150 1301 2202
rect 1301 2150 1311 2202
rect 1335 2150 1365 2202
rect 1365 2150 1377 2202
rect 1377 2150 1391 2202
rect 1415 2150 1429 2202
rect 1429 2150 1441 2202
rect 1441 2150 1471 2202
rect 1495 2150 1505 2202
rect 1505 2150 1551 2202
rect 1255 2148 1311 2150
rect 1335 2148 1391 2150
rect 1415 2148 1471 2150
rect 1495 2148 1551 2150
rect 2957 2202 3013 2204
rect 3037 2202 3093 2204
rect 3117 2202 3173 2204
rect 3197 2202 3253 2204
rect 2957 2150 3003 2202
rect 3003 2150 3013 2202
rect 3037 2150 3067 2202
rect 3067 2150 3079 2202
rect 3079 2150 3093 2202
rect 3117 2150 3131 2202
rect 3131 2150 3143 2202
rect 3143 2150 3173 2202
rect 3197 2150 3207 2202
rect 3207 2150 3253 2202
rect 2957 2148 3013 2150
rect 3037 2148 3093 2150
rect 3117 2148 3173 2150
rect 3197 2148 3253 2150
rect 4659 2202 4715 2204
rect 4739 2202 4795 2204
rect 4819 2202 4875 2204
rect 4899 2202 4955 2204
rect 4659 2150 4705 2202
rect 4705 2150 4715 2202
rect 4739 2150 4769 2202
rect 4769 2150 4781 2202
rect 4781 2150 4795 2202
rect 4819 2150 4833 2202
rect 4833 2150 4845 2202
rect 4845 2150 4875 2202
rect 4899 2150 4909 2202
rect 4909 2150 4955 2202
rect 4659 2148 4715 2150
rect 4739 2148 4795 2150
rect 4819 2148 4875 2150
rect 4899 2148 4955 2150
rect 6361 2202 6417 2204
rect 6441 2202 6497 2204
rect 6521 2202 6577 2204
rect 6601 2202 6657 2204
rect 6361 2150 6407 2202
rect 6407 2150 6417 2202
rect 6441 2150 6471 2202
rect 6471 2150 6483 2202
rect 6483 2150 6497 2202
rect 6521 2150 6535 2202
rect 6535 2150 6547 2202
rect 6547 2150 6577 2202
rect 6601 2150 6611 2202
rect 6611 2150 6657 2202
rect 6361 2148 6417 2150
rect 6441 2148 6497 2150
rect 6521 2148 6577 2150
rect 6601 2148 6657 2150
rect 2106 1658 2162 1660
rect 2186 1658 2242 1660
rect 2266 1658 2322 1660
rect 2346 1658 2402 1660
rect 2106 1606 2152 1658
rect 2152 1606 2162 1658
rect 2186 1606 2216 1658
rect 2216 1606 2228 1658
rect 2228 1606 2242 1658
rect 2266 1606 2280 1658
rect 2280 1606 2292 1658
rect 2292 1606 2322 1658
rect 2346 1606 2356 1658
rect 2356 1606 2402 1658
rect 2106 1604 2162 1606
rect 2186 1604 2242 1606
rect 2266 1604 2322 1606
rect 2346 1604 2402 1606
rect 3808 1658 3864 1660
rect 3888 1658 3944 1660
rect 3968 1658 4024 1660
rect 4048 1658 4104 1660
rect 3808 1606 3854 1658
rect 3854 1606 3864 1658
rect 3888 1606 3918 1658
rect 3918 1606 3930 1658
rect 3930 1606 3944 1658
rect 3968 1606 3982 1658
rect 3982 1606 3994 1658
rect 3994 1606 4024 1658
rect 4048 1606 4058 1658
rect 4058 1606 4104 1658
rect 3808 1604 3864 1606
rect 3888 1604 3944 1606
rect 3968 1604 4024 1606
rect 4048 1604 4104 1606
rect 5510 1658 5566 1660
rect 5590 1658 5646 1660
rect 5670 1658 5726 1660
rect 5750 1658 5806 1660
rect 5510 1606 5556 1658
rect 5556 1606 5566 1658
rect 5590 1606 5620 1658
rect 5620 1606 5632 1658
rect 5632 1606 5646 1658
rect 5670 1606 5684 1658
rect 5684 1606 5696 1658
rect 5696 1606 5726 1658
rect 5750 1606 5760 1658
rect 5760 1606 5806 1658
rect 5510 1604 5566 1606
rect 5590 1604 5646 1606
rect 5670 1604 5726 1606
rect 5750 1604 5806 1606
rect 7212 1658 7268 1660
rect 7292 1658 7348 1660
rect 7372 1658 7428 1660
rect 7452 1658 7508 1660
rect 7212 1606 7258 1658
rect 7258 1606 7268 1658
rect 7292 1606 7322 1658
rect 7322 1606 7334 1658
rect 7334 1606 7348 1658
rect 7372 1606 7386 1658
rect 7386 1606 7398 1658
rect 7398 1606 7428 1658
rect 7452 1606 7462 1658
rect 7462 1606 7508 1658
rect 7212 1604 7268 1606
rect 7292 1604 7348 1606
rect 7372 1604 7428 1606
rect 7452 1604 7508 1606
rect 1255 1114 1311 1116
rect 1335 1114 1391 1116
rect 1415 1114 1471 1116
rect 1495 1114 1551 1116
rect 1255 1062 1301 1114
rect 1301 1062 1311 1114
rect 1335 1062 1365 1114
rect 1365 1062 1377 1114
rect 1377 1062 1391 1114
rect 1415 1062 1429 1114
rect 1429 1062 1441 1114
rect 1441 1062 1471 1114
rect 1495 1062 1505 1114
rect 1505 1062 1551 1114
rect 1255 1060 1311 1062
rect 1335 1060 1391 1062
rect 1415 1060 1471 1062
rect 1495 1060 1551 1062
rect 2957 1114 3013 1116
rect 3037 1114 3093 1116
rect 3117 1114 3173 1116
rect 3197 1114 3253 1116
rect 2957 1062 3003 1114
rect 3003 1062 3013 1114
rect 3037 1062 3067 1114
rect 3067 1062 3079 1114
rect 3079 1062 3093 1114
rect 3117 1062 3131 1114
rect 3131 1062 3143 1114
rect 3143 1062 3173 1114
rect 3197 1062 3207 1114
rect 3207 1062 3253 1114
rect 2957 1060 3013 1062
rect 3037 1060 3093 1062
rect 3117 1060 3173 1062
rect 3197 1060 3253 1062
rect 4659 1114 4715 1116
rect 4739 1114 4795 1116
rect 4819 1114 4875 1116
rect 4899 1114 4955 1116
rect 4659 1062 4705 1114
rect 4705 1062 4715 1114
rect 4739 1062 4769 1114
rect 4769 1062 4781 1114
rect 4781 1062 4795 1114
rect 4819 1062 4833 1114
rect 4833 1062 4845 1114
rect 4845 1062 4875 1114
rect 4899 1062 4909 1114
rect 4909 1062 4955 1114
rect 4659 1060 4715 1062
rect 4739 1060 4795 1062
rect 4819 1060 4875 1062
rect 4899 1060 4955 1062
rect 6361 1114 6417 1116
rect 6441 1114 6497 1116
rect 6521 1114 6577 1116
rect 6601 1114 6657 1116
rect 6361 1062 6407 1114
rect 6407 1062 6417 1114
rect 6441 1062 6471 1114
rect 6471 1062 6483 1114
rect 6483 1062 6497 1114
rect 6521 1062 6535 1114
rect 6535 1062 6547 1114
rect 6547 1062 6577 1114
rect 6601 1062 6611 1114
rect 6611 1062 6657 1114
rect 6361 1060 6417 1062
rect 6441 1060 6497 1062
rect 6521 1060 6577 1062
rect 6601 1060 6657 1062
rect 2106 570 2162 572
rect 2186 570 2242 572
rect 2266 570 2322 572
rect 2346 570 2402 572
rect 2106 518 2152 570
rect 2152 518 2162 570
rect 2186 518 2216 570
rect 2216 518 2228 570
rect 2228 518 2242 570
rect 2266 518 2280 570
rect 2280 518 2292 570
rect 2292 518 2322 570
rect 2346 518 2356 570
rect 2356 518 2402 570
rect 2106 516 2162 518
rect 2186 516 2242 518
rect 2266 516 2322 518
rect 2346 516 2402 518
rect 3808 570 3864 572
rect 3888 570 3944 572
rect 3968 570 4024 572
rect 4048 570 4104 572
rect 3808 518 3854 570
rect 3854 518 3864 570
rect 3888 518 3918 570
rect 3918 518 3930 570
rect 3930 518 3944 570
rect 3968 518 3982 570
rect 3982 518 3994 570
rect 3994 518 4024 570
rect 4048 518 4058 570
rect 4058 518 4104 570
rect 3808 516 3864 518
rect 3888 516 3944 518
rect 3968 516 4024 518
rect 4048 516 4104 518
rect 5510 570 5566 572
rect 5590 570 5646 572
rect 5670 570 5726 572
rect 5750 570 5806 572
rect 5510 518 5556 570
rect 5556 518 5566 570
rect 5590 518 5620 570
rect 5620 518 5632 570
rect 5632 518 5646 570
rect 5670 518 5684 570
rect 5684 518 5696 570
rect 5696 518 5726 570
rect 5750 518 5760 570
rect 5760 518 5806 570
rect 5510 516 5566 518
rect 5590 516 5646 518
rect 5670 516 5726 518
rect 5750 516 5806 518
rect 7212 570 7268 572
rect 7292 570 7348 572
rect 7372 570 7428 572
rect 7452 570 7508 572
rect 7212 518 7258 570
rect 7258 518 7268 570
rect 7292 518 7322 570
rect 7322 518 7334 570
rect 7334 518 7348 570
rect 7372 518 7386 570
rect 7386 518 7398 570
rect 7398 518 7428 570
rect 7452 518 7462 570
rect 7462 518 7508 570
rect 7212 516 7268 518
rect 7292 516 7348 518
rect 7372 516 7428 518
rect 7452 516 7508 518
<< metal3 >>
rect 2096 7104 2412 7105
rect 2096 7040 2102 7104
rect 2166 7040 2182 7104
rect 2246 7040 2262 7104
rect 2326 7040 2342 7104
rect 2406 7040 2412 7104
rect 2096 7039 2412 7040
rect 3798 7104 4114 7105
rect 3798 7040 3804 7104
rect 3868 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4114 7104
rect 3798 7039 4114 7040
rect 5500 7104 5816 7105
rect 5500 7040 5506 7104
rect 5570 7040 5586 7104
rect 5650 7040 5666 7104
rect 5730 7040 5746 7104
rect 5810 7040 5816 7104
rect 5500 7039 5816 7040
rect 7202 7104 7518 7105
rect 7202 7040 7208 7104
rect 7272 7040 7288 7104
rect 7352 7040 7368 7104
rect 7432 7040 7448 7104
rect 7512 7040 7518 7104
rect 7202 7039 7518 7040
rect 1245 6560 1561 6561
rect 1245 6496 1251 6560
rect 1315 6496 1331 6560
rect 1395 6496 1411 6560
rect 1475 6496 1491 6560
rect 1555 6496 1561 6560
rect 1245 6495 1561 6496
rect 2947 6560 3263 6561
rect 2947 6496 2953 6560
rect 3017 6496 3033 6560
rect 3097 6496 3113 6560
rect 3177 6496 3193 6560
rect 3257 6496 3263 6560
rect 2947 6495 3263 6496
rect 4649 6560 4965 6561
rect 4649 6496 4655 6560
rect 4719 6496 4735 6560
rect 4799 6496 4815 6560
rect 4879 6496 4895 6560
rect 4959 6496 4965 6560
rect 4649 6495 4965 6496
rect 6351 6560 6667 6561
rect 6351 6496 6357 6560
rect 6421 6496 6437 6560
rect 6501 6496 6517 6560
rect 6581 6496 6597 6560
rect 6661 6496 6667 6560
rect 6351 6495 6667 6496
rect 2096 6016 2412 6017
rect 2096 5952 2102 6016
rect 2166 5952 2182 6016
rect 2246 5952 2262 6016
rect 2326 5952 2342 6016
rect 2406 5952 2412 6016
rect 2096 5951 2412 5952
rect 3798 6016 4114 6017
rect 3798 5952 3804 6016
rect 3868 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4114 6016
rect 3798 5951 4114 5952
rect 5500 6016 5816 6017
rect 5500 5952 5506 6016
rect 5570 5952 5586 6016
rect 5650 5952 5666 6016
rect 5730 5952 5746 6016
rect 5810 5952 5816 6016
rect 5500 5951 5816 5952
rect 7202 6016 7518 6017
rect 7202 5952 7208 6016
rect 7272 5952 7288 6016
rect 7352 5952 7368 6016
rect 7432 5952 7448 6016
rect 7512 5952 7518 6016
rect 7202 5951 7518 5952
rect 1245 5472 1561 5473
rect 1245 5408 1251 5472
rect 1315 5408 1331 5472
rect 1395 5408 1411 5472
rect 1475 5408 1491 5472
rect 1555 5408 1561 5472
rect 1245 5407 1561 5408
rect 2947 5472 3263 5473
rect 2947 5408 2953 5472
rect 3017 5408 3033 5472
rect 3097 5408 3113 5472
rect 3177 5408 3193 5472
rect 3257 5408 3263 5472
rect 2947 5407 3263 5408
rect 4649 5472 4965 5473
rect 4649 5408 4655 5472
rect 4719 5408 4735 5472
rect 4799 5408 4815 5472
rect 4879 5408 4895 5472
rect 4959 5408 4965 5472
rect 4649 5407 4965 5408
rect 6351 5472 6667 5473
rect 6351 5408 6357 5472
rect 6421 5408 6437 5472
rect 6501 5408 6517 5472
rect 6581 5408 6597 5472
rect 6661 5408 6667 5472
rect 6351 5407 6667 5408
rect 2096 4928 2412 4929
rect 2096 4864 2102 4928
rect 2166 4864 2182 4928
rect 2246 4864 2262 4928
rect 2326 4864 2342 4928
rect 2406 4864 2412 4928
rect 2096 4863 2412 4864
rect 3798 4928 4114 4929
rect 3798 4864 3804 4928
rect 3868 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4114 4928
rect 3798 4863 4114 4864
rect 5500 4928 5816 4929
rect 5500 4864 5506 4928
rect 5570 4864 5586 4928
rect 5650 4864 5666 4928
rect 5730 4864 5746 4928
rect 5810 4864 5816 4928
rect 5500 4863 5816 4864
rect 7202 4928 7518 4929
rect 7202 4864 7208 4928
rect 7272 4864 7288 4928
rect 7352 4864 7368 4928
rect 7432 4864 7448 4928
rect 7512 4864 7518 4928
rect 7202 4863 7518 4864
rect 1245 4384 1561 4385
rect 1245 4320 1251 4384
rect 1315 4320 1331 4384
rect 1395 4320 1411 4384
rect 1475 4320 1491 4384
rect 1555 4320 1561 4384
rect 1245 4319 1561 4320
rect 2947 4384 3263 4385
rect 2947 4320 2953 4384
rect 3017 4320 3033 4384
rect 3097 4320 3113 4384
rect 3177 4320 3193 4384
rect 3257 4320 3263 4384
rect 2947 4319 3263 4320
rect 4649 4384 4965 4385
rect 4649 4320 4655 4384
rect 4719 4320 4735 4384
rect 4799 4320 4815 4384
rect 4879 4320 4895 4384
rect 4959 4320 4965 4384
rect 4649 4319 4965 4320
rect 6351 4384 6667 4385
rect 6351 4320 6357 4384
rect 6421 4320 6437 4384
rect 6501 4320 6517 4384
rect 6581 4320 6597 4384
rect 6661 4320 6667 4384
rect 6351 4319 6667 4320
rect 2096 3840 2412 3841
rect 2096 3776 2102 3840
rect 2166 3776 2182 3840
rect 2246 3776 2262 3840
rect 2326 3776 2342 3840
rect 2406 3776 2412 3840
rect 2096 3775 2412 3776
rect 3798 3840 4114 3841
rect 3798 3776 3804 3840
rect 3868 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4114 3840
rect 3798 3775 4114 3776
rect 5500 3840 5816 3841
rect 5500 3776 5506 3840
rect 5570 3776 5586 3840
rect 5650 3776 5666 3840
rect 5730 3776 5746 3840
rect 5810 3776 5816 3840
rect 5500 3775 5816 3776
rect 7202 3840 7518 3841
rect 7202 3776 7208 3840
rect 7272 3776 7288 3840
rect 7352 3776 7368 3840
rect 7432 3776 7448 3840
rect 7512 3776 7518 3840
rect 7202 3775 7518 3776
rect 1245 3296 1561 3297
rect 1245 3232 1251 3296
rect 1315 3232 1331 3296
rect 1395 3232 1411 3296
rect 1475 3232 1491 3296
rect 1555 3232 1561 3296
rect 1245 3231 1561 3232
rect 2947 3296 3263 3297
rect 2947 3232 2953 3296
rect 3017 3232 3033 3296
rect 3097 3232 3113 3296
rect 3177 3232 3193 3296
rect 3257 3232 3263 3296
rect 2947 3231 3263 3232
rect 4649 3296 4965 3297
rect 4649 3232 4655 3296
rect 4719 3232 4735 3296
rect 4799 3232 4815 3296
rect 4879 3232 4895 3296
rect 4959 3232 4965 3296
rect 4649 3231 4965 3232
rect 6351 3296 6667 3297
rect 6351 3232 6357 3296
rect 6421 3232 6437 3296
rect 6501 3232 6517 3296
rect 6581 3232 6597 3296
rect 6661 3232 6667 3296
rect 6351 3231 6667 3232
rect 2096 2752 2412 2753
rect 2096 2688 2102 2752
rect 2166 2688 2182 2752
rect 2246 2688 2262 2752
rect 2326 2688 2342 2752
rect 2406 2688 2412 2752
rect 2096 2687 2412 2688
rect 3798 2752 4114 2753
rect 3798 2688 3804 2752
rect 3868 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4114 2752
rect 3798 2687 4114 2688
rect 5500 2752 5816 2753
rect 5500 2688 5506 2752
rect 5570 2688 5586 2752
rect 5650 2688 5666 2752
rect 5730 2688 5746 2752
rect 5810 2688 5816 2752
rect 5500 2687 5816 2688
rect 7202 2752 7518 2753
rect 7202 2688 7208 2752
rect 7272 2688 7288 2752
rect 7352 2688 7368 2752
rect 7432 2688 7448 2752
rect 7512 2688 7518 2752
rect 7202 2687 7518 2688
rect 1245 2208 1561 2209
rect 1245 2144 1251 2208
rect 1315 2144 1331 2208
rect 1395 2144 1411 2208
rect 1475 2144 1491 2208
rect 1555 2144 1561 2208
rect 1245 2143 1561 2144
rect 2947 2208 3263 2209
rect 2947 2144 2953 2208
rect 3017 2144 3033 2208
rect 3097 2144 3113 2208
rect 3177 2144 3193 2208
rect 3257 2144 3263 2208
rect 2947 2143 3263 2144
rect 4649 2208 4965 2209
rect 4649 2144 4655 2208
rect 4719 2144 4735 2208
rect 4799 2144 4815 2208
rect 4879 2144 4895 2208
rect 4959 2144 4965 2208
rect 4649 2143 4965 2144
rect 6351 2208 6667 2209
rect 6351 2144 6357 2208
rect 6421 2144 6437 2208
rect 6501 2144 6517 2208
rect 6581 2144 6597 2208
rect 6661 2144 6667 2208
rect 6351 2143 6667 2144
rect 2096 1664 2412 1665
rect 2096 1600 2102 1664
rect 2166 1600 2182 1664
rect 2246 1600 2262 1664
rect 2326 1600 2342 1664
rect 2406 1600 2412 1664
rect 2096 1599 2412 1600
rect 3798 1664 4114 1665
rect 3798 1600 3804 1664
rect 3868 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4114 1664
rect 3798 1599 4114 1600
rect 5500 1664 5816 1665
rect 5500 1600 5506 1664
rect 5570 1600 5586 1664
rect 5650 1600 5666 1664
rect 5730 1600 5746 1664
rect 5810 1600 5816 1664
rect 5500 1599 5816 1600
rect 7202 1664 7518 1665
rect 7202 1600 7208 1664
rect 7272 1600 7288 1664
rect 7352 1600 7368 1664
rect 7432 1600 7448 1664
rect 7512 1600 7518 1664
rect 7202 1599 7518 1600
rect 1245 1120 1561 1121
rect 1245 1056 1251 1120
rect 1315 1056 1331 1120
rect 1395 1056 1411 1120
rect 1475 1056 1491 1120
rect 1555 1056 1561 1120
rect 1245 1055 1561 1056
rect 2947 1120 3263 1121
rect 2947 1056 2953 1120
rect 3017 1056 3033 1120
rect 3097 1056 3113 1120
rect 3177 1056 3193 1120
rect 3257 1056 3263 1120
rect 2947 1055 3263 1056
rect 4649 1120 4965 1121
rect 4649 1056 4655 1120
rect 4719 1056 4735 1120
rect 4799 1056 4815 1120
rect 4879 1056 4895 1120
rect 4959 1056 4965 1120
rect 4649 1055 4965 1056
rect 6351 1120 6667 1121
rect 6351 1056 6357 1120
rect 6421 1056 6437 1120
rect 6501 1056 6517 1120
rect 6581 1056 6597 1120
rect 6661 1056 6667 1120
rect 6351 1055 6667 1056
rect 2096 576 2412 577
rect 2096 512 2102 576
rect 2166 512 2182 576
rect 2246 512 2262 576
rect 2326 512 2342 576
rect 2406 512 2412 576
rect 2096 511 2412 512
rect 3798 576 4114 577
rect 3798 512 3804 576
rect 3868 512 3884 576
rect 3948 512 3964 576
rect 4028 512 4044 576
rect 4108 512 4114 576
rect 3798 511 4114 512
rect 5500 576 5816 577
rect 5500 512 5506 576
rect 5570 512 5586 576
rect 5650 512 5666 576
rect 5730 512 5746 576
rect 5810 512 5816 576
rect 5500 511 5816 512
rect 7202 576 7518 577
rect 7202 512 7208 576
rect 7272 512 7288 576
rect 7352 512 7368 576
rect 7432 512 7448 576
rect 7512 512 7518 576
rect 7202 511 7518 512
<< via3 >>
rect 2102 7100 2166 7104
rect 2102 7044 2106 7100
rect 2106 7044 2162 7100
rect 2162 7044 2166 7100
rect 2102 7040 2166 7044
rect 2182 7100 2246 7104
rect 2182 7044 2186 7100
rect 2186 7044 2242 7100
rect 2242 7044 2246 7100
rect 2182 7040 2246 7044
rect 2262 7100 2326 7104
rect 2262 7044 2266 7100
rect 2266 7044 2322 7100
rect 2322 7044 2326 7100
rect 2262 7040 2326 7044
rect 2342 7100 2406 7104
rect 2342 7044 2346 7100
rect 2346 7044 2402 7100
rect 2402 7044 2406 7100
rect 2342 7040 2406 7044
rect 3804 7100 3868 7104
rect 3804 7044 3808 7100
rect 3808 7044 3864 7100
rect 3864 7044 3868 7100
rect 3804 7040 3868 7044
rect 3884 7100 3948 7104
rect 3884 7044 3888 7100
rect 3888 7044 3944 7100
rect 3944 7044 3948 7100
rect 3884 7040 3948 7044
rect 3964 7100 4028 7104
rect 3964 7044 3968 7100
rect 3968 7044 4024 7100
rect 4024 7044 4028 7100
rect 3964 7040 4028 7044
rect 4044 7100 4108 7104
rect 4044 7044 4048 7100
rect 4048 7044 4104 7100
rect 4104 7044 4108 7100
rect 4044 7040 4108 7044
rect 5506 7100 5570 7104
rect 5506 7044 5510 7100
rect 5510 7044 5566 7100
rect 5566 7044 5570 7100
rect 5506 7040 5570 7044
rect 5586 7100 5650 7104
rect 5586 7044 5590 7100
rect 5590 7044 5646 7100
rect 5646 7044 5650 7100
rect 5586 7040 5650 7044
rect 5666 7100 5730 7104
rect 5666 7044 5670 7100
rect 5670 7044 5726 7100
rect 5726 7044 5730 7100
rect 5666 7040 5730 7044
rect 5746 7100 5810 7104
rect 5746 7044 5750 7100
rect 5750 7044 5806 7100
rect 5806 7044 5810 7100
rect 5746 7040 5810 7044
rect 7208 7100 7272 7104
rect 7208 7044 7212 7100
rect 7212 7044 7268 7100
rect 7268 7044 7272 7100
rect 7208 7040 7272 7044
rect 7288 7100 7352 7104
rect 7288 7044 7292 7100
rect 7292 7044 7348 7100
rect 7348 7044 7352 7100
rect 7288 7040 7352 7044
rect 7368 7100 7432 7104
rect 7368 7044 7372 7100
rect 7372 7044 7428 7100
rect 7428 7044 7432 7100
rect 7368 7040 7432 7044
rect 7448 7100 7512 7104
rect 7448 7044 7452 7100
rect 7452 7044 7508 7100
rect 7508 7044 7512 7100
rect 7448 7040 7512 7044
rect 1251 6556 1315 6560
rect 1251 6500 1255 6556
rect 1255 6500 1311 6556
rect 1311 6500 1315 6556
rect 1251 6496 1315 6500
rect 1331 6556 1395 6560
rect 1331 6500 1335 6556
rect 1335 6500 1391 6556
rect 1391 6500 1395 6556
rect 1331 6496 1395 6500
rect 1411 6556 1475 6560
rect 1411 6500 1415 6556
rect 1415 6500 1471 6556
rect 1471 6500 1475 6556
rect 1411 6496 1475 6500
rect 1491 6556 1555 6560
rect 1491 6500 1495 6556
rect 1495 6500 1551 6556
rect 1551 6500 1555 6556
rect 1491 6496 1555 6500
rect 2953 6556 3017 6560
rect 2953 6500 2957 6556
rect 2957 6500 3013 6556
rect 3013 6500 3017 6556
rect 2953 6496 3017 6500
rect 3033 6556 3097 6560
rect 3033 6500 3037 6556
rect 3037 6500 3093 6556
rect 3093 6500 3097 6556
rect 3033 6496 3097 6500
rect 3113 6556 3177 6560
rect 3113 6500 3117 6556
rect 3117 6500 3173 6556
rect 3173 6500 3177 6556
rect 3113 6496 3177 6500
rect 3193 6556 3257 6560
rect 3193 6500 3197 6556
rect 3197 6500 3253 6556
rect 3253 6500 3257 6556
rect 3193 6496 3257 6500
rect 4655 6556 4719 6560
rect 4655 6500 4659 6556
rect 4659 6500 4715 6556
rect 4715 6500 4719 6556
rect 4655 6496 4719 6500
rect 4735 6556 4799 6560
rect 4735 6500 4739 6556
rect 4739 6500 4795 6556
rect 4795 6500 4799 6556
rect 4735 6496 4799 6500
rect 4815 6556 4879 6560
rect 4815 6500 4819 6556
rect 4819 6500 4875 6556
rect 4875 6500 4879 6556
rect 4815 6496 4879 6500
rect 4895 6556 4959 6560
rect 4895 6500 4899 6556
rect 4899 6500 4955 6556
rect 4955 6500 4959 6556
rect 4895 6496 4959 6500
rect 6357 6556 6421 6560
rect 6357 6500 6361 6556
rect 6361 6500 6417 6556
rect 6417 6500 6421 6556
rect 6357 6496 6421 6500
rect 6437 6556 6501 6560
rect 6437 6500 6441 6556
rect 6441 6500 6497 6556
rect 6497 6500 6501 6556
rect 6437 6496 6501 6500
rect 6517 6556 6581 6560
rect 6517 6500 6521 6556
rect 6521 6500 6577 6556
rect 6577 6500 6581 6556
rect 6517 6496 6581 6500
rect 6597 6556 6661 6560
rect 6597 6500 6601 6556
rect 6601 6500 6657 6556
rect 6657 6500 6661 6556
rect 6597 6496 6661 6500
rect 2102 6012 2166 6016
rect 2102 5956 2106 6012
rect 2106 5956 2162 6012
rect 2162 5956 2166 6012
rect 2102 5952 2166 5956
rect 2182 6012 2246 6016
rect 2182 5956 2186 6012
rect 2186 5956 2242 6012
rect 2242 5956 2246 6012
rect 2182 5952 2246 5956
rect 2262 6012 2326 6016
rect 2262 5956 2266 6012
rect 2266 5956 2322 6012
rect 2322 5956 2326 6012
rect 2262 5952 2326 5956
rect 2342 6012 2406 6016
rect 2342 5956 2346 6012
rect 2346 5956 2402 6012
rect 2402 5956 2406 6012
rect 2342 5952 2406 5956
rect 3804 6012 3868 6016
rect 3804 5956 3808 6012
rect 3808 5956 3864 6012
rect 3864 5956 3868 6012
rect 3804 5952 3868 5956
rect 3884 6012 3948 6016
rect 3884 5956 3888 6012
rect 3888 5956 3944 6012
rect 3944 5956 3948 6012
rect 3884 5952 3948 5956
rect 3964 6012 4028 6016
rect 3964 5956 3968 6012
rect 3968 5956 4024 6012
rect 4024 5956 4028 6012
rect 3964 5952 4028 5956
rect 4044 6012 4108 6016
rect 4044 5956 4048 6012
rect 4048 5956 4104 6012
rect 4104 5956 4108 6012
rect 4044 5952 4108 5956
rect 5506 6012 5570 6016
rect 5506 5956 5510 6012
rect 5510 5956 5566 6012
rect 5566 5956 5570 6012
rect 5506 5952 5570 5956
rect 5586 6012 5650 6016
rect 5586 5956 5590 6012
rect 5590 5956 5646 6012
rect 5646 5956 5650 6012
rect 5586 5952 5650 5956
rect 5666 6012 5730 6016
rect 5666 5956 5670 6012
rect 5670 5956 5726 6012
rect 5726 5956 5730 6012
rect 5666 5952 5730 5956
rect 5746 6012 5810 6016
rect 5746 5956 5750 6012
rect 5750 5956 5806 6012
rect 5806 5956 5810 6012
rect 5746 5952 5810 5956
rect 7208 6012 7272 6016
rect 7208 5956 7212 6012
rect 7212 5956 7268 6012
rect 7268 5956 7272 6012
rect 7208 5952 7272 5956
rect 7288 6012 7352 6016
rect 7288 5956 7292 6012
rect 7292 5956 7348 6012
rect 7348 5956 7352 6012
rect 7288 5952 7352 5956
rect 7368 6012 7432 6016
rect 7368 5956 7372 6012
rect 7372 5956 7428 6012
rect 7428 5956 7432 6012
rect 7368 5952 7432 5956
rect 7448 6012 7512 6016
rect 7448 5956 7452 6012
rect 7452 5956 7508 6012
rect 7508 5956 7512 6012
rect 7448 5952 7512 5956
rect 1251 5468 1315 5472
rect 1251 5412 1255 5468
rect 1255 5412 1311 5468
rect 1311 5412 1315 5468
rect 1251 5408 1315 5412
rect 1331 5468 1395 5472
rect 1331 5412 1335 5468
rect 1335 5412 1391 5468
rect 1391 5412 1395 5468
rect 1331 5408 1395 5412
rect 1411 5468 1475 5472
rect 1411 5412 1415 5468
rect 1415 5412 1471 5468
rect 1471 5412 1475 5468
rect 1411 5408 1475 5412
rect 1491 5468 1555 5472
rect 1491 5412 1495 5468
rect 1495 5412 1551 5468
rect 1551 5412 1555 5468
rect 1491 5408 1555 5412
rect 2953 5468 3017 5472
rect 2953 5412 2957 5468
rect 2957 5412 3013 5468
rect 3013 5412 3017 5468
rect 2953 5408 3017 5412
rect 3033 5468 3097 5472
rect 3033 5412 3037 5468
rect 3037 5412 3093 5468
rect 3093 5412 3097 5468
rect 3033 5408 3097 5412
rect 3113 5468 3177 5472
rect 3113 5412 3117 5468
rect 3117 5412 3173 5468
rect 3173 5412 3177 5468
rect 3113 5408 3177 5412
rect 3193 5468 3257 5472
rect 3193 5412 3197 5468
rect 3197 5412 3253 5468
rect 3253 5412 3257 5468
rect 3193 5408 3257 5412
rect 4655 5468 4719 5472
rect 4655 5412 4659 5468
rect 4659 5412 4715 5468
rect 4715 5412 4719 5468
rect 4655 5408 4719 5412
rect 4735 5468 4799 5472
rect 4735 5412 4739 5468
rect 4739 5412 4795 5468
rect 4795 5412 4799 5468
rect 4735 5408 4799 5412
rect 4815 5468 4879 5472
rect 4815 5412 4819 5468
rect 4819 5412 4875 5468
rect 4875 5412 4879 5468
rect 4815 5408 4879 5412
rect 4895 5468 4959 5472
rect 4895 5412 4899 5468
rect 4899 5412 4955 5468
rect 4955 5412 4959 5468
rect 4895 5408 4959 5412
rect 6357 5468 6421 5472
rect 6357 5412 6361 5468
rect 6361 5412 6417 5468
rect 6417 5412 6421 5468
rect 6357 5408 6421 5412
rect 6437 5468 6501 5472
rect 6437 5412 6441 5468
rect 6441 5412 6497 5468
rect 6497 5412 6501 5468
rect 6437 5408 6501 5412
rect 6517 5468 6581 5472
rect 6517 5412 6521 5468
rect 6521 5412 6577 5468
rect 6577 5412 6581 5468
rect 6517 5408 6581 5412
rect 6597 5468 6661 5472
rect 6597 5412 6601 5468
rect 6601 5412 6657 5468
rect 6657 5412 6661 5468
rect 6597 5408 6661 5412
rect 2102 4924 2166 4928
rect 2102 4868 2106 4924
rect 2106 4868 2162 4924
rect 2162 4868 2166 4924
rect 2102 4864 2166 4868
rect 2182 4924 2246 4928
rect 2182 4868 2186 4924
rect 2186 4868 2242 4924
rect 2242 4868 2246 4924
rect 2182 4864 2246 4868
rect 2262 4924 2326 4928
rect 2262 4868 2266 4924
rect 2266 4868 2322 4924
rect 2322 4868 2326 4924
rect 2262 4864 2326 4868
rect 2342 4924 2406 4928
rect 2342 4868 2346 4924
rect 2346 4868 2402 4924
rect 2402 4868 2406 4924
rect 2342 4864 2406 4868
rect 3804 4924 3868 4928
rect 3804 4868 3808 4924
rect 3808 4868 3864 4924
rect 3864 4868 3868 4924
rect 3804 4864 3868 4868
rect 3884 4924 3948 4928
rect 3884 4868 3888 4924
rect 3888 4868 3944 4924
rect 3944 4868 3948 4924
rect 3884 4864 3948 4868
rect 3964 4924 4028 4928
rect 3964 4868 3968 4924
rect 3968 4868 4024 4924
rect 4024 4868 4028 4924
rect 3964 4864 4028 4868
rect 4044 4924 4108 4928
rect 4044 4868 4048 4924
rect 4048 4868 4104 4924
rect 4104 4868 4108 4924
rect 4044 4864 4108 4868
rect 5506 4924 5570 4928
rect 5506 4868 5510 4924
rect 5510 4868 5566 4924
rect 5566 4868 5570 4924
rect 5506 4864 5570 4868
rect 5586 4924 5650 4928
rect 5586 4868 5590 4924
rect 5590 4868 5646 4924
rect 5646 4868 5650 4924
rect 5586 4864 5650 4868
rect 5666 4924 5730 4928
rect 5666 4868 5670 4924
rect 5670 4868 5726 4924
rect 5726 4868 5730 4924
rect 5666 4864 5730 4868
rect 5746 4924 5810 4928
rect 5746 4868 5750 4924
rect 5750 4868 5806 4924
rect 5806 4868 5810 4924
rect 5746 4864 5810 4868
rect 7208 4924 7272 4928
rect 7208 4868 7212 4924
rect 7212 4868 7268 4924
rect 7268 4868 7272 4924
rect 7208 4864 7272 4868
rect 7288 4924 7352 4928
rect 7288 4868 7292 4924
rect 7292 4868 7348 4924
rect 7348 4868 7352 4924
rect 7288 4864 7352 4868
rect 7368 4924 7432 4928
rect 7368 4868 7372 4924
rect 7372 4868 7428 4924
rect 7428 4868 7432 4924
rect 7368 4864 7432 4868
rect 7448 4924 7512 4928
rect 7448 4868 7452 4924
rect 7452 4868 7508 4924
rect 7508 4868 7512 4924
rect 7448 4864 7512 4868
rect 1251 4380 1315 4384
rect 1251 4324 1255 4380
rect 1255 4324 1311 4380
rect 1311 4324 1315 4380
rect 1251 4320 1315 4324
rect 1331 4380 1395 4384
rect 1331 4324 1335 4380
rect 1335 4324 1391 4380
rect 1391 4324 1395 4380
rect 1331 4320 1395 4324
rect 1411 4380 1475 4384
rect 1411 4324 1415 4380
rect 1415 4324 1471 4380
rect 1471 4324 1475 4380
rect 1411 4320 1475 4324
rect 1491 4380 1555 4384
rect 1491 4324 1495 4380
rect 1495 4324 1551 4380
rect 1551 4324 1555 4380
rect 1491 4320 1555 4324
rect 2953 4380 3017 4384
rect 2953 4324 2957 4380
rect 2957 4324 3013 4380
rect 3013 4324 3017 4380
rect 2953 4320 3017 4324
rect 3033 4380 3097 4384
rect 3033 4324 3037 4380
rect 3037 4324 3093 4380
rect 3093 4324 3097 4380
rect 3033 4320 3097 4324
rect 3113 4380 3177 4384
rect 3113 4324 3117 4380
rect 3117 4324 3173 4380
rect 3173 4324 3177 4380
rect 3113 4320 3177 4324
rect 3193 4380 3257 4384
rect 3193 4324 3197 4380
rect 3197 4324 3253 4380
rect 3253 4324 3257 4380
rect 3193 4320 3257 4324
rect 4655 4380 4719 4384
rect 4655 4324 4659 4380
rect 4659 4324 4715 4380
rect 4715 4324 4719 4380
rect 4655 4320 4719 4324
rect 4735 4380 4799 4384
rect 4735 4324 4739 4380
rect 4739 4324 4795 4380
rect 4795 4324 4799 4380
rect 4735 4320 4799 4324
rect 4815 4380 4879 4384
rect 4815 4324 4819 4380
rect 4819 4324 4875 4380
rect 4875 4324 4879 4380
rect 4815 4320 4879 4324
rect 4895 4380 4959 4384
rect 4895 4324 4899 4380
rect 4899 4324 4955 4380
rect 4955 4324 4959 4380
rect 4895 4320 4959 4324
rect 6357 4380 6421 4384
rect 6357 4324 6361 4380
rect 6361 4324 6417 4380
rect 6417 4324 6421 4380
rect 6357 4320 6421 4324
rect 6437 4380 6501 4384
rect 6437 4324 6441 4380
rect 6441 4324 6497 4380
rect 6497 4324 6501 4380
rect 6437 4320 6501 4324
rect 6517 4380 6581 4384
rect 6517 4324 6521 4380
rect 6521 4324 6577 4380
rect 6577 4324 6581 4380
rect 6517 4320 6581 4324
rect 6597 4380 6661 4384
rect 6597 4324 6601 4380
rect 6601 4324 6657 4380
rect 6657 4324 6661 4380
rect 6597 4320 6661 4324
rect 2102 3836 2166 3840
rect 2102 3780 2106 3836
rect 2106 3780 2162 3836
rect 2162 3780 2166 3836
rect 2102 3776 2166 3780
rect 2182 3836 2246 3840
rect 2182 3780 2186 3836
rect 2186 3780 2242 3836
rect 2242 3780 2246 3836
rect 2182 3776 2246 3780
rect 2262 3836 2326 3840
rect 2262 3780 2266 3836
rect 2266 3780 2322 3836
rect 2322 3780 2326 3836
rect 2262 3776 2326 3780
rect 2342 3836 2406 3840
rect 2342 3780 2346 3836
rect 2346 3780 2402 3836
rect 2402 3780 2406 3836
rect 2342 3776 2406 3780
rect 3804 3836 3868 3840
rect 3804 3780 3808 3836
rect 3808 3780 3864 3836
rect 3864 3780 3868 3836
rect 3804 3776 3868 3780
rect 3884 3836 3948 3840
rect 3884 3780 3888 3836
rect 3888 3780 3944 3836
rect 3944 3780 3948 3836
rect 3884 3776 3948 3780
rect 3964 3836 4028 3840
rect 3964 3780 3968 3836
rect 3968 3780 4024 3836
rect 4024 3780 4028 3836
rect 3964 3776 4028 3780
rect 4044 3836 4108 3840
rect 4044 3780 4048 3836
rect 4048 3780 4104 3836
rect 4104 3780 4108 3836
rect 4044 3776 4108 3780
rect 5506 3836 5570 3840
rect 5506 3780 5510 3836
rect 5510 3780 5566 3836
rect 5566 3780 5570 3836
rect 5506 3776 5570 3780
rect 5586 3836 5650 3840
rect 5586 3780 5590 3836
rect 5590 3780 5646 3836
rect 5646 3780 5650 3836
rect 5586 3776 5650 3780
rect 5666 3836 5730 3840
rect 5666 3780 5670 3836
rect 5670 3780 5726 3836
rect 5726 3780 5730 3836
rect 5666 3776 5730 3780
rect 5746 3836 5810 3840
rect 5746 3780 5750 3836
rect 5750 3780 5806 3836
rect 5806 3780 5810 3836
rect 5746 3776 5810 3780
rect 7208 3836 7272 3840
rect 7208 3780 7212 3836
rect 7212 3780 7268 3836
rect 7268 3780 7272 3836
rect 7208 3776 7272 3780
rect 7288 3836 7352 3840
rect 7288 3780 7292 3836
rect 7292 3780 7348 3836
rect 7348 3780 7352 3836
rect 7288 3776 7352 3780
rect 7368 3836 7432 3840
rect 7368 3780 7372 3836
rect 7372 3780 7428 3836
rect 7428 3780 7432 3836
rect 7368 3776 7432 3780
rect 7448 3836 7512 3840
rect 7448 3780 7452 3836
rect 7452 3780 7508 3836
rect 7508 3780 7512 3836
rect 7448 3776 7512 3780
rect 1251 3292 1315 3296
rect 1251 3236 1255 3292
rect 1255 3236 1311 3292
rect 1311 3236 1315 3292
rect 1251 3232 1315 3236
rect 1331 3292 1395 3296
rect 1331 3236 1335 3292
rect 1335 3236 1391 3292
rect 1391 3236 1395 3292
rect 1331 3232 1395 3236
rect 1411 3292 1475 3296
rect 1411 3236 1415 3292
rect 1415 3236 1471 3292
rect 1471 3236 1475 3292
rect 1411 3232 1475 3236
rect 1491 3292 1555 3296
rect 1491 3236 1495 3292
rect 1495 3236 1551 3292
rect 1551 3236 1555 3292
rect 1491 3232 1555 3236
rect 2953 3292 3017 3296
rect 2953 3236 2957 3292
rect 2957 3236 3013 3292
rect 3013 3236 3017 3292
rect 2953 3232 3017 3236
rect 3033 3292 3097 3296
rect 3033 3236 3037 3292
rect 3037 3236 3093 3292
rect 3093 3236 3097 3292
rect 3033 3232 3097 3236
rect 3113 3292 3177 3296
rect 3113 3236 3117 3292
rect 3117 3236 3173 3292
rect 3173 3236 3177 3292
rect 3113 3232 3177 3236
rect 3193 3292 3257 3296
rect 3193 3236 3197 3292
rect 3197 3236 3253 3292
rect 3253 3236 3257 3292
rect 3193 3232 3257 3236
rect 4655 3292 4719 3296
rect 4655 3236 4659 3292
rect 4659 3236 4715 3292
rect 4715 3236 4719 3292
rect 4655 3232 4719 3236
rect 4735 3292 4799 3296
rect 4735 3236 4739 3292
rect 4739 3236 4795 3292
rect 4795 3236 4799 3292
rect 4735 3232 4799 3236
rect 4815 3292 4879 3296
rect 4815 3236 4819 3292
rect 4819 3236 4875 3292
rect 4875 3236 4879 3292
rect 4815 3232 4879 3236
rect 4895 3292 4959 3296
rect 4895 3236 4899 3292
rect 4899 3236 4955 3292
rect 4955 3236 4959 3292
rect 4895 3232 4959 3236
rect 6357 3292 6421 3296
rect 6357 3236 6361 3292
rect 6361 3236 6417 3292
rect 6417 3236 6421 3292
rect 6357 3232 6421 3236
rect 6437 3292 6501 3296
rect 6437 3236 6441 3292
rect 6441 3236 6497 3292
rect 6497 3236 6501 3292
rect 6437 3232 6501 3236
rect 6517 3292 6581 3296
rect 6517 3236 6521 3292
rect 6521 3236 6577 3292
rect 6577 3236 6581 3292
rect 6517 3232 6581 3236
rect 6597 3292 6661 3296
rect 6597 3236 6601 3292
rect 6601 3236 6657 3292
rect 6657 3236 6661 3292
rect 6597 3232 6661 3236
rect 2102 2748 2166 2752
rect 2102 2692 2106 2748
rect 2106 2692 2162 2748
rect 2162 2692 2166 2748
rect 2102 2688 2166 2692
rect 2182 2748 2246 2752
rect 2182 2692 2186 2748
rect 2186 2692 2242 2748
rect 2242 2692 2246 2748
rect 2182 2688 2246 2692
rect 2262 2748 2326 2752
rect 2262 2692 2266 2748
rect 2266 2692 2322 2748
rect 2322 2692 2326 2748
rect 2262 2688 2326 2692
rect 2342 2748 2406 2752
rect 2342 2692 2346 2748
rect 2346 2692 2402 2748
rect 2402 2692 2406 2748
rect 2342 2688 2406 2692
rect 3804 2748 3868 2752
rect 3804 2692 3808 2748
rect 3808 2692 3864 2748
rect 3864 2692 3868 2748
rect 3804 2688 3868 2692
rect 3884 2748 3948 2752
rect 3884 2692 3888 2748
rect 3888 2692 3944 2748
rect 3944 2692 3948 2748
rect 3884 2688 3948 2692
rect 3964 2748 4028 2752
rect 3964 2692 3968 2748
rect 3968 2692 4024 2748
rect 4024 2692 4028 2748
rect 3964 2688 4028 2692
rect 4044 2748 4108 2752
rect 4044 2692 4048 2748
rect 4048 2692 4104 2748
rect 4104 2692 4108 2748
rect 4044 2688 4108 2692
rect 5506 2748 5570 2752
rect 5506 2692 5510 2748
rect 5510 2692 5566 2748
rect 5566 2692 5570 2748
rect 5506 2688 5570 2692
rect 5586 2748 5650 2752
rect 5586 2692 5590 2748
rect 5590 2692 5646 2748
rect 5646 2692 5650 2748
rect 5586 2688 5650 2692
rect 5666 2748 5730 2752
rect 5666 2692 5670 2748
rect 5670 2692 5726 2748
rect 5726 2692 5730 2748
rect 5666 2688 5730 2692
rect 5746 2748 5810 2752
rect 5746 2692 5750 2748
rect 5750 2692 5806 2748
rect 5806 2692 5810 2748
rect 5746 2688 5810 2692
rect 7208 2748 7272 2752
rect 7208 2692 7212 2748
rect 7212 2692 7268 2748
rect 7268 2692 7272 2748
rect 7208 2688 7272 2692
rect 7288 2748 7352 2752
rect 7288 2692 7292 2748
rect 7292 2692 7348 2748
rect 7348 2692 7352 2748
rect 7288 2688 7352 2692
rect 7368 2748 7432 2752
rect 7368 2692 7372 2748
rect 7372 2692 7428 2748
rect 7428 2692 7432 2748
rect 7368 2688 7432 2692
rect 7448 2748 7512 2752
rect 7448 2692 7452 2748
rect 7452 2692 7508 2748
rect 7508 2692 7512 2748
rect 7448 2688 7512 2692
rect 1251 2204 1315 2208
rect 1251 2148 1255 2204
rect 1255 2148 1311 2204
rect 1311 2148 1315 2204
rect 1251 2144 1315 2148
rect 1331 2204 1395 2208
rect 1331 2148 1335 2204
rect 1335 2148 1391 2204
rect 1391 2148 1395 2204
rect 1331 2144 1395 2148
rect 1411 2204 1475 2208
rect 1411 2148 1415 2204
rect 1415 2148 1471 2204
rect 1471 2148 1475 2204
rect 1411 2144 1475 2148
rect 1491 2204 1555 2208
rect 1491 2148 1495 2204
rect 1495 2148 1551 2204
rect 1551 2148 1555 2204
rect 1491 2144 1555 2148
rect 2953 2204 3017 2208
rect 2953 2148 2957 2204
rect 2957 2148 3013 2204
rect 3013 2148 3017 2204
rect 2953 2144 3017 2148
rect 3033 2204 3097 2208
rect 3033 2148 3037 2204
rect 3037 2148 3093 2204
rect 3093 2148 3097 2204
rect 3033 2144 3097 2148
rect 3113 2204 3177 2208
rect 3113 2148 3117 2204
rect 3117 2148 3173 2204
rect 3173 2148 3177 2204
rect 3113 2144 3177 2148
rect 3193 2204 3257 2208
rect 3193 2148 3197 2204
rect 3197 2148 3253 2204
rect 3253 2148 3257 2204
rect 3193 2144 3257 2148
rect 4655 2204 4719 2208
rect 4655 2148 4659 2204
rect 4659 2148 4715 2204
rect 4715 2148 4719 2204
rect 4655 2144 4719 2148
rect 4735 2204 4799 2208
rect 4735 2148 4739 2204
rect 4739 2148 4795 2204
rect 4795 2148 4799 2204
rect 4735 2144 4799 2148
rect 4815 2204 4879 2208
rect 4815 2148 4819 2204
rect 4819 2148 4875 2204
rect 4875 2148 4879 2204
rect 4815 2144 4879 2148
rect 4895 2204 4959 2208
rect 4895 2148 4899 2204
rect 4899 2148 4955 2204
rect 4955 2148 4959 2204
rect 4895 2144 4959 2148
rect 6357 2204 6421 2208
rect 6357 2148 6361 2204
rect 6361 2148 6417 2204
rect 6417 2148 6421 2204
rect 6357 2144 6421 2148
rect 6437 2204 6501 2208
rect 6437 2148 6441 2204
rect 6441 2148 6497 2204
rect 6497 2148 6501 2204
rect 6437 2144 6501 2148
rect 6517 2204 6581 2208
rect 6517 2148 6521 2204
rect 6521 2148 6577 2204
rect 6577 2148 6581 2204
rect 6517 2144 6581 2148
rect 6597 2204 6661 2208
rect 6597 2148 6601 2204
rect 6601 2148 6657 2204
rect 6657 2148 6661 2204
rect 6597 2144 6661 2148
rect 2102 1660 2166 1664
rect 2102 1604 2106 1660
rect 2106 1604 2162 1660
rect 2162 1604 2166 1660
rect 2102 1600 2166 1604
rect 2182 1660 2246 1664
rect 2182 1604 2186 1660
rect 2186 1604 2242 1660
rect 2242 1604 2246 1660
rect 2182 1600 2246 1604
rect 2262 1660 2326 1664
rect 2262 1604 2266 1660
rect 2266 1604 2322 1660
rect 2322 1604 2326 1660
rect 2262 1600 2326 1604
rect 2342 1660 2406 1664
rect 2342 1604 2346 1660
rect 2346 1604 2402 1660
rect 2402 1604 2406 1660
rect 2342 1600 2406 1604
rect 3804 1660 3868 1664
rect 3804 1604 3808 1660
rect 3808 1604 3864 1660
rect 3864 1604 3868 1660
rect 3804 1600 3868 1604
rect 3884 1660 3948 1664
rect 3884 1604 3888 1660
rect 3888 1604 3944 1660
rect 3944 1604 3948 1660
rect 3884 1600 3948 1604
rect 3964 1660 4028 1664
rect 3964 1604 3968 1660
rect 3968 1604 4024 1660
rect 4024 1604 4028 1660
rect 3964 1600 4028 1604
rect 4044 1660 4108 1664
rect 4044 1604 4048 1660
rect 4048 1604 4104 1660
rect 4104 1604 4108 1660
rect 4044 1600 4108 1604
rect 5506 1660 5570 1664
rect 5506 1604 5510 1660
rect 5510 1604 5566 1660
rect 5566 1604 5570 1660
rect 5506 1600 5570 1604
rect 5586 1660 5650 1664
rect 5586 1604 5590 1660
rect 5590 1604 5646 1660
rect 5646 1604 5650 1660
rect 5586 1600 5650 1604
rect 5666 1660 5730 1664
rect 5666 1604 5670 1660
rect 5670 1604 5726 1660
rect 5726 1604 5730 1660
rect 5666 1600 5730 1604
rect 5746 1660 5810 1664
rect 5746 1604 5750 1660
rect 5750 1604 5806 1660
rect 5806 1604 5810 1660
rect 5746 1600 5810 1604
rect 7208 1660 7272 1664
rect 7208 1604 7212 1660
rect 7212 1604 7268 1660
rect 7268 1604 7272 1660
rect 7208 1600 7272 1604
rect 7288 1660 7352 1664
rect 7288 1604 7292 1660
rect 7292 1604 7348 1660
rect 7348 1604 7352 1660
rect 7288 1600 7352 1604
rect 7368 1660 7432 1664
rect 7368 1604 7372 1660
rect 7372 1604 7428 1660
rect 7428 1604 7432 1660
rect 7368 1600 7432 1604
rect 7448 1660 7512 1664
rect 7448 1604 7452 1660
rect 7452 1604 7508 1660
rect 7508 1604 7512 1660
rect 7448 1600 7512 1604
rect 1251 1116 1315 1120
rect 1251 1060 1255 1116
rect 1255 1060 1311 1116
rect 1311 1060 1315 1116
rect 1251 1056 1315 1060
rect 1331 1116 1395 1120
rect 1331 1060 1335 1116
rect 1335 1060 1391 1116
rect 1391 1060 1395 1116
rect 1331 1056 1395 1060
rect 1411 1116 1475 1120
rect 1411 1060 1415 1116
rect 1415 1060 1471 1116
rect 1471 1060 1475 1116
rect 1411 1056 1475 1060
rect 1491 1116 1555 1120
rect 1491 1060 1495 1116
rect 1495 1060 1551 1116
rect 1551 1060 1555 1116
rect 1491 1056 1555 1060
rect 2953 1116 3017 1120
rect 2953 1060 2957 1116
rect 2957 1060 3013 1116
rect 3013 1060 3017 1116
rect 2953 1056 3017 1060
rect 3033 1116 3097 1120
rect 3033 1060 3037 1116
rect 3037 1060 3093 1116
rect 3093 1060 3097 1116
rect 3033 1056 3097 1060
rect 3113 1116 3177 1120
rect 3113 1060 3117 1116
rect 3117 1060 3173 1116
rect 3173 1060 3177 1116
rect 3113 1056 3177 1060
rect 3193 1116 3257 1120
rect 3193 1060 3197 1116
rect 3197 1060 3253 1116
rect 3253 1060 3257 1116
rect 3193 1056 3257 1060
rect 4655 1116 4719 1120
rect 4655 1060 4659 1116
rect 4659 1060 4715 1116
rect 4715 1060 4719 1116
rect 4655 1056 4719 1060
rect 4735 1116 4799 1120
rect 4735 1060 4739 1116
rect 4739 1060 4795 1116
rect 4795 1060 4799 1116
rect 4735 1056 4799 1060
rect 4815 1116 4879 1120
rect 4815 1060 4819 1116
rect 4819 1060 4875 1116
rect 4875 1060 4879 1116
rect 4815 1056 4879 1060
rect 4895 1116 4959 1120
rect 4895 1060 4899 1116
rect 4899 1060 4955 1116
rect 4955 1060 4959 1116
rect 4895 1056 4959 1060
rect 6357 1116 6421 1120
rect 6357 1060 6361 1116
rect 6361 1060 6417 1116
rect 6417 1060 6421 1116
rect 6357 1056 6421 1060
rect 6437 1116 6501 1120
rect 6437 1060 6441 1116
rect 6441 1060 6497 1116
rect 6497 1060 6501 1116
rect 6437 1056 6501 1060
rect 6517 1116 6581 1120
rect 6517 1060 6521 1116
rect 6521 1060 6577 1116
rect 6577 1060 6581 1116
rect 6517 1056 6581 1060
rect 6597 1116 6661 1120
rect 6597 1060 6601 1116
rect 6601 1060 6657 1116
rect 6657 1060 6661 1116
rect 6597 1056 6661 1060
rect 2102 572 2166 576
rect 2102 516 2106 572
rect 2106 516 2162 572
rect 2162 516 2166 572
rect 2102 512 2166 516
rect 2182 572 2246 576
rect 2182 516 2186 572
rect 2186 516 2242 572
rect 2242 516 2246 572
rect 2182 512 2246 516
rect 2262 572 2326 576
rect 2262 516 2266 572
rect 2266 516 2322 572
rect 2322 516 2326 572
rect 2262 512 2326 516
rect 2342 572 2406 576
rect 2342 516 2346 572
rect 2346 516 2402 572
rect 2402 516 2406 572
rect 2342 512 2406 516
rect 3804 572 3868 576
rect 3804 516 3808 572
rect 3808 516 3864 572
rect 3864 516 3868 572
rect 3804 512 3868 516
rect 3884 572 3948 576
rect 3884 516 3888 572
rect 3888 516 3944 572
rect 3944 516 3948 572
rect 3884 512 3948 516
rect 3964 572 4028 576
rect 3964 516 3968 572
rect 3968 516 4024 572
rect 4024 516 4028 572
rect 3964 512 4028 516
rect 4044 572 4108 576
rect 4044 516 4048 572
rect 4048 516 4104 572
rect 4104 516 4108 572
rect 4044 512 4108 516
rect 5506 572 5570 576
rect 5506 516 5510 572
rect 5510 516 5566 572
rect 5566 516 5570 572
rect 5506 512 5570 516
rect 5586 572 5650 576
rect 5586 516 5590 572
rect 5590 516 5646 572
rect 5646 516 5650 572
rect 5586 512 5650 516
rect 5666 572 5730 576
rect 5666 516 5670 572
rect 5670 516 5726 572
rect 5726 516 5730 572
rect 5666 512 5730 516
rect 5746 572 5810 576
rect 5746 516 5750 572
rect 5750 516 5806 572
rect 5806 516 5810 572
rect 5746 512 5810 516
rect 7208 572 7272 576
rect 7208 516 7212 572
rect 7212 516 7268 572
rect 7268 516 7272 572
rect 7208 512 7272 516
rect 7288 572 7352 576
rect 7288 516 7292 572
rect 7292 516 7348 572
rect 7348 516 7352 572
rect 7288 512 7352 516
rect 7368 572 7432 576
rect 7368 516 7372 572
rect 7372 516 7428 572
rect 7428 516 7432 572
rect 7368 512 7432 516
rect 7448 572 7512 576
rect 7448 516 7452 572
rect 7452 516 7508 572
rect 7508 516 7512 572
rect 7448 512 7512 516
<< metal4 >>
rect 1243 6560 1563 7120
rect 1243 6496 1251 6560
rect 1315 6496 1331 6560
rect 1395 6496 1411 6560
rect 1475 6496 1491 6560
rect 1555 6496 1563 6560
rect 1243 5472 1563 6496
rect 1243 5408 1251 5472
rect 1315 5408 1331 5472
rect 1395 5408 1411 5472
rect 1475 5408 1491 5472
rect 1555 5408 1563 5472
rect 1243 4384 1563 5408
rect 1243 4320 1251 4384
rect 1315 4320 1331 4384
rect 1395 4320 1411 4384
rect 1475 4320 1491 4384
rect 1555 4320 1563 4384
rect 1243 3296 1563 4320
rect 1243 3232 1251 3296
rect 1315 3232 1331 3296
rect 1395 3232 1411 3296
rect 1475 3232 1491 3296
rect 1555 3232 1563 3296
rect 1243 2208 1563 3232
rect 1243 2144 1251 2208
rect 1315 2144 1331 2208
rect 1395 2144 1411 2208
rect 1475 2144 1491 2208
rect 1555 2144 1563 2208
rect 1243 1120 1563 2144
rect 1243 1056 1251 1120
rect 1315 1056 1331 1120
rect 1395 1056 1411 1120
rect 1475 1056 1491 1120
rect 1555 1056 1563 1120
rect 1243 496 1563 1056
rect 2094 7104 2414 7120
rect 2094 7040 2102 7104
rect 2166 7040 2182 7104
rect 2246 7040 2262 7104
rect 2326 7040 2342 7104
rect 2406 7040 2414 7104
rect 2094 6016 2414 7040
rect 2094 5952 2102 6016
rect 2166 5952 2182 6016
rect 2246 5952 2262 6016
rect 2326 5952 2342 6016
rect 2406 5952 2414 6016
rect 2094 4928 2414 5952
rect 2094 4864 2102 4928
rect 2166 4864 2182 4928
rect 2246 4864 2262 4928
rect 2326 4864 2342 4928
rect 2406 4864 2414 4928
rect 2094 3840 2414 4864
rect 2094 3776 2102 3840
rect 2166 3776 2182 3840
rect 2246 3776 2262 3840
rect 2326 3776 2342 3840
rect 2406 3776 2414 3840
rect 2094 2752 2414 3776
rect 2094 2688 2102 2752
rect 2166 2688 2182 2752
rect 2246 2688 2262 2752
rect 2326 2688 2342 2752
rect 2406 2688 2414 2752
rect 2094 1664 2414 2688
rect 2094 1600 2102 1664
rect 2166 1600 2182 1664
rect 2246 1600 2262 1664
rect 2326 1600 2342 1664
rect 2406 1600 2414 1664
rect 2094 576 2414 1600
rect 2094 512 2102 576
rect 2166 512 2182 576
rect 2246 512 2262 576
rect 2326 512 2342 576
rect 2406 512 2414 576
rect 2094 496 2414 512
rect 2945 6560 3265 7120
rect 2945 6496 2953 6560
rect 3017 6496 3033 6560
rect 3097 6496 3113 6560
rect 3177 6496 3193 6560
rect 3257 6496 3265 6560
rect 2945 5472 3265 6496
rect 2945 5408 2953 5472
rect 3017 5408 3033 5472
rect 3097 5408 3113 5472
rect 3177 5408 3193 5472
rect 3257 5408 3265 5472
rect 2945 4384 3265 5408
rect 2945 4320 2953 4384
rect 3017 4320 3033 4384
rect 3097 4320 3113 4384
rect 3177 4320 3193 4384
rect 3257 4320 3265 4384
rect 2945 3296 3265 4320
rect 2945 3232 2953 3296
rect 3017 3232 3033 3296
rect 3097 3232 3113 3296
rect 3177 3232 3193 3296
rect 3257 3232 3265 3296
rect 2945 2208 3265 3232
rect 2945 2144 2953 2208
rect 3017 2144 3033 2208
rect 3097 2144 3113 2208
rect 3177 2144 3193 2208
rect 3257 2144 3265 2208
rect 2945 1120 3265 2144
rect 2945 1056 2953 1120
rect 3017 1056 3033 1120
rect 3097 1056 3113 1120
rect 3177 1056 3193 1120
rect 3257 1056 3265 1120
rect 2945 496 3265 1056
rect 3796 7104 4116 7120
rect 3796 7040 3804 7104
rect 3868 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4116 7104
rect 3796 6016 4116 7040
rect 3796 5952 3804 6016
rect 3868 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4116 6016
rect 3796 4928 4116 5952
rect 3796 4864 3804 4928
rect 3868 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4116 4928
rect 3796 3840 4116 4864
rect 3796 3776 3804 3840
rect 3868 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4116 3840
rect 3796 2752 4116 3776
rect 3796 2688 3804 2752
rect 3868 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4116 2752
rect 3796 1664 4116 2688
rect 3796 1600 3804 1664
rect 3868 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4116 1664
rect 3796 576 4116 1600
rect 3796 512 3804 576
rect 3868 512 3884 576
rect 3948 512 3964 576
rect 4028 512 4044 576
rect 4108 512 4116 576
rect 3796 496 4116 512
rect 4647 6560 4967 7120
rect 4647 6496 4655 6560
rect 4719 6496 4735 6560
rect 4799 6496 4815 6560
rect 4879 6496 4895 6560
rect 4959 6496 4967 6560
rect 4647 5472 4967 6496
rect 4647 5408 4655 5472
rect 4719 5408 4735 5472
rect 4799 5408 4815 5472
rect 4879 5408 4895 5472
rect 4959 5408 4967 5472
rect 4647 4384 4967 5408
rect 4647 4320 4655 4384
rect 4719 4320 4735 4384
rect 4799 4320 4815 4384
rect 4879 4320 4895 4384
rect 4959 4320 4967 4384
rect 4647 3296 4967 4320
rect 4647 3232 4655 3296
rect 4719 3232 4735 3296
rect 4799 3232 4815 3296
rect 4879 3232 4895 3296
rect 4959 3232 4967 3296
rect 4647 2208 4967 3232
rect 4647 2144 4655 2208
rect 4719 2144 4735 2208
rect 4799 2144 4815 2208
rect 4879 2144 4895 2208
rect 4959 2144 4967 2208
rect 4647 1120 4967 2144
rect 4647 1056 4655 1120
rect 4719 1056 4735 1120
rect 4799 1056 4815 1120
rect 4879 1056 4895 1120
rect 4959 1056 4967 1120
rect 4647 496 4967 1056
rect 5498 7104 5818 7120
rect 5498 7040 5506 7104
rect 5570 7040 5586 7104
rect 5650 7040 5666 7104
rect 5730 7040 5746 7104
rect 5810 7040 5818 7104
rect 5498 6016 5818 7040
rect 5498 5952 5506 6016
rect 5570 5952 5586 6016
rect 5650 5952 5666 6016
rect 5730 5952 5746 6016
rect 5810 5952 5818 6016
rect 5498 4928 5818 5952
rect 5498 4864 5506 4928
rect 5570 4864 5586 4928
rect 5650 4864 5666 4928
rect 5730 4864 5746 4928
rect 5810 4864 5818 4928
rect 5498 3840 5818 4864
rect 5498 3776 5506 3840
rect 5570 3776 5586 3840
rect 5650 3776 5666 3840
rect 5730 3776 5746 3840
rect 5810 3776 5818 3840
rect 5498 2752 5818 3776
rect 5498 2688 5506 2752
rect 5570 2688 5586 2752
rect 5650 2688 5666 2752
rect 5730 2688 5746 2752
rect 5810 2688 5818 2752
rect 5498 1664 5818 2688
rect 5498 1600 5506 1664
rect 5570 1600 5586 1664
rect 5650 1600 5666 1664
rect 5730 1600 5746 1664
rect 5810 1600 5818 1664
rect 5498 576 5818 1600
rect 5498 512 5506 576
rect 5570 512 5586 576
rect 5650 512 5666 576
rect 5730 512 5746 576
rect 5810 512 5818 576
rect 5498 496 5818 512
rect 6349 6560 6669 7120
rect 6349 6496 6357 6560
rect 6421 6496 6437 6560
rect 6501 6496 6517 6560
rect 6581 6496 6597 6560
rect 6661 6496 6669 6560
rect 6349 5472 6669 6496
rect 6349 5408 6357 5472
rect 6421 5408 6437 5472
rect 6501 5408 6517 5472
rect 6581 5408 6597 5472
rect 6661 5408 6669 5472
rect 6349 4384 6669 5408
rect 6349 4320 6357 4384
rect 6421 4320 6437 4384
rect 6501 4320 6517 4384
rect 6581 4320 6597 4384
rect 6661 4320 6669 4384
rect 6349 3296 6669 4320
rect 6349 3232 6357 3296
rect 6421 3232 6437 3296
rect 6501 3232 6517 3296
rect 6581 3232 6597 3296
rect 6661 3232 6669 3296
rect 6349 2208 6669 3232
rect 6349 2144 6357 2208
rect 6421 2144 6437 2208
rect 6501 2144 6517 2208
rect 6581 2144 6597 2208
rect 6661 2144 6669 2208
rect 6349 1120 6669 2144
rect 6349 1056 6357 1120
rect 6421 1056 6437 1120
rect 6501 1056 6517 1120
rect 6581 1056 6597 1120
rect 6661 1056 6669 1120
rect 6349 496 6669 1056
rect 7200 7104 7520 7120
rect 7200 7040 7208 7104
rect 7272 7040 7288 7104
rect 7352 7040 7368 7104
rect 7432 7040 7448 7104
rect 7512 7040 7520 7104
rect 7200 6016 7520 7040
rect 7200 5952 7208 6016
rect 7272 5952 7288 6016
rect 7352 5952 7368 6016
rect 7432 5952 7448 6016
rect 7512 5952 7520 6016
rect 7200 4928 7520 5952
rect 7200 4864 7208 4928
rect 7272 4864 7288 4928
rect 7352 4864 7368 4928
rect 7432 4864 7448 4928
rect 7512 4864 7520 4928
rect 7200 3840 7520 4864
rect 7200 3776 7208 3840
rect 7272 3776 7288 3840
rect 7352 3776 7368 3840
rect 7432 3776 7448 3840
rect 7512 3776 7520 3840
rect 7200 2752 7520 3776
rect 7200 2688 7208 2752
rect 7272 2688 7288 2752
rect 7352 2688 7368 2752
rect 7432 2688 7448 2752
rect 7512 2688 7520 2752
rect 7200 1664 7520 2688
rect 7200 1600 7208 1664
rect 7272 1600 7288 1664
rect 7352 1600 7368 1664
rect 7432 1600 7448 1664
rect 7512 1600 7520 1664
rect 7200 576 7520 1600
rect 7200 512 7208 576
rect 7272 512 7288 576
rect 7352 512 7368 576
rect 7432 512 7448 576
rect 7512 512 7520 576
rect 7200 496 7520 512
use sky130_fd_sc_hd__inv_2  _1_
timestamp 0
transform 1 0 3956 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2_
timestamp 0
transform -1 0 3772 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _3_
timestamp 0
transform -1 0 3864 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _4_
timestamp 0
transform -1 0 2944 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _5_
timestamp 0
transform -1 0 4508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _6_
timestamp 0
transform 1 0 3772 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _7_
timestamp 0
transform -1 0 5520 0 1 4896
box -38 -48 1970 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69
timestamp 0
transform 1 0 6900 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_69
timestamp 0
transform 1 0 6900 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_65
timestamp 0
transform 1 0 6532 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 0
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_65
timestamp 0
transform 1 0 6532 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 0
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_65
timestamp 0
transform 1 0 6532 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_69
timestamp 0
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 0
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 0
transform 1 0 5520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_66
timestamp 0
transform 1 0 6624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_70
timestamp 0
transform 1 0 6992 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 0
transform 1 0 1932 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_19
timestamp 0
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_69
timestamp 0
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 0
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_36
timestamp 0
transform 1 0 3864 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_43
timestamp 0
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_47
timestamp 0
transform 1 0 4876 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_56
timestamp 0
transform 1 0 5704 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_68
timestamp 0
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_27
timestamp 0
transform 1 0 3036 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_29
timestamp 0
transform 1 0 3220 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_41
timestamp 0
transform 1 0 4324 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 0
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 0
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_65
timestamp 0
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 5704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 7360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 7360 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 7360 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 7360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 7360 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 7360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 7360 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 0
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 0
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 0
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 0
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 0
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 0
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 0
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 0
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 0
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 0
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 0
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 0
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 0
transform 1 0 3128 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 0
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
<< labels >>
rlabel metal2 s 4036 7072 4036 7072 4 VGND
rlabel metal1 s 3956 6528 3956 6528 4 VPWR
rlabel metal1 s 2806 5848 2806 5848 4 _0_
rlabel metal1 s 3818 5814 3818 5814 4 clk
rlabel metal1 s 4232 5814 4232 5814 4 f0.d
rlabel metal1 s 3358 5746 3358 5746 4 f0.q
rlabel metal1 s 4692 5202 4692 5202 4 f1.d
rlabel metal2 s 3726 5542 3726 5542 4 f1.q
rlabel metal1 s 6946 6834 6946 6834 4 n_rst
rlabel metal1 s 5343 5814 5343 5814 4 net1
rlabel metal1 s 4738 6222 4738 6222 4 net2
rlabel metal2 s 2937 7684 2937 7684 4 out_i
rlabel metal1 s 2024 5814 2024 5814 4 out_q
flabel metal4 s 7200 496 7520 7120 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5498 496 5818 7120 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3796 496 4116 7120 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2094 496 2414 7120 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6349 496 6669 7120 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4647 496 4967 7120 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2945 496 3265 7120 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1243 496 1563 7120 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 4894 7600 4950 8000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 6826 7600 6882 8000 0 FreeSans 280 90 0 0 n_rst
port 4 nsew
flabel metal2 s 2962 7600 3018 8000 0 FreeSans 280 90 0 0 out_i
port 5 nsew
flabel metal2 s 1030 7600 1086 8000 0 FreeSans 280 90 0 0 out_q
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 8000 8000
string GDS_END 144964
string GDS_FILE ../gds/quadrature_divider.gds
string GDS_START 68118
<< end >>
