magic
tech sky130A
magscale 1 2
timestamp 1716495612
<< pwell >>
rect -1083 -1210 1083 1210
<< nmos >>
rect -887 -1000 -487 1000
rect -429 -1000 -29 1000
rect 29 -1000 429 1000
rect 487 -1000 887 1000
<< ndiff >>
rect -945 988 -887 1000
rect -945 -988 -933 988
rect -899 -988 -887 988
rect -945 -1000 -887 -988
rect -487 988 -429 1000
rect -487 -988 -475 988
rect -441 -988 -429 988
rect -487 -1000 -429 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 429 988 487 1000
rect 429 -988 441 988
rect 475 -988 487 988
rect 429 -1000 487 -988
rect 887 988 945 1000
rect 887 -988 899 988
rect 933 -988 945 988
rect 887 -1000 945 -988
<< ndiffc >>
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
<< psubdiff >>
rect -1047 1140 -951 1174
rect 951 1140 1047 1174
rect -1047 1078 -1013 1140
rect 1013 1078 1047 1140
rect -1047 -1140 -1013 -1078
rect 1013 -1140 1047 -1078
rect -1047 -1174 -951 -1140
rect 951 -1174 1047 -1140
<< psubdiffcont >>
rect -951 1140 951 1174
rect -1047 -1078 -1013 1078
rect 1013 -1078 1047 1078
rect -951 -1174 951 -1140
<< poly >>
rect -887 1072 -487 1088
rect -887 1038 -871 1072
rect -503 1038 -487 1072
rect -887 1000 -487 1038
rect -429 1072 -29 1088
rect -429 1038 -413 1072
rect -45 1038 -29 1072
rect -429 1000 -29 1038
rect 29 1072 429 1088
rect 29 1038 45 1072
rect 413 1038 429 1072
rect 29 1000 429 1038
rect 487 1072 887 1088
rect 487 1038 503 1072
rect 871 1038 887 1072
rect 487 1000 887 1038
rect -887 -1038 -487 -1000
rect -887 -1072 -871 -1038
rect -503 -1072 -487 -1038
rect -887 -1088 -487 -1072
rect -429 -1038 -29 -1000
rect -429 -1072 -413 -1038
rect -45 -1072 -29 -1038
rect -429 -1088 -29 -1072
rect 29 -1038 429 -1000
rect 29 -1072 45 -1038
rect 413 -1072 429 -1038
rect 29 -1088 429 -1072
rect 487 -1038 887 -1000
rect 487 -1072 503 -1038
rect 871 -1072 887 -1038
rect 487 -1088 887 -1072
<< polycont >>
rect -871 1038 -503 1072
rect -413 1038 -45 1072
rect 45 1038 413 1072
rect 503 1038 871 1072
rect -871 -1072 -503 -1038
rect -413 -1072 -45 -1038
rect 45 -1072 413 -1038
rect 503 -1072 871 -1038
<< locali >>
rect -1047 1140 -951 1174
rect 951 1140 1047 1174
rect -1047 1078 -1013 1140
rect 1013 1078 1047 1140
rect -887 1038 -871 1072
rect -503 1038 -487 1072
rect -429 1038 -413 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 413 1038 429 1072
rect 487 1038 503 1072
rect 871 1038 887 1072
rect -933 988 -899 1004
rect -933 -1004 -899 -988
rect -475 988 -441 1004
rect -475 -1004 -441 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 441 988 475 1004
rect 441 -1004 475 -988
rect 899 988 933 1004
rect 899 -1004 933 -988
rect -887 -1072 -871 -1038
rect -503 -1072 -487 -1038
rect -429 -1072 -413 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 413 -1072 429 -1038
rect 487 -1072 503 -1038
rect 871 -1072 887 -1038
rect -1047 -1140 -1013 -1078
rect 1013 -1140 1047 -1078
rect -1047 -1174 -951 -1140
rect 951 -1174 1047 -1140
<< viali >>
rect -871 1038 -503 1072
rect -413 1038 -45 1072
rect 45 1038 413 1072
rect 503 1038 871 1072
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
rect -871 -1072 -503 -1038
rect -413 -1072 -45 -1038
rect 45 -1072 413 -1038
rect 503 -1072 871 -1038
<< metal1 >>
rect -883 1072 -491 1078
rect -883 1038 -871 1072
rect -503 1038 -491 1072
rect -883 1032 -491 1038
rect -425 1072 -33 1078
rect -425 1038 -413 1072
rect -45 1038 -33 1072
rect -425 1032 -33 1038
rect 33 1072 425 1078
rect 33 1038 45 1072
rect 413 1038 425 1072
rect 33 1032 425 1038
rect 491 1072 883 1078
rect 491 1038 503 1072
rect 871 1038 883 1072
rect 491 1032 883 1038
rect -939 988 -893 1000
rect -939 -988 -933 988
rect -899 -988 -893 988
rect -939 -1000 -893 -988
rect -481 988 -435 1000
rect -481 -988 -475 988
rect -441 -988 -435 988
rect -481 -1000 -435 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 435 988 481 1000
rect 435 -988 441 988
rect 475 -988 481 988
rect 435 -1000 481 -988
rect 893 988 939 1000
rect 893 -988 899 988
rect 933 -988 939 988
rect 893 -1000 939 -988
rect -883 -1038 -491 -1032
rect -883 -1072 -871 -1038
rect -503 -1072 -491 -1038
rect -883 -1078 -491 -1072
rect -425 -1038 -33 -1032
rect -425 -1072 -413 -1038
rect -45 -1072 -33 -1038
rect -425 -1078 -33 -1072
rect 33 -1038 425 -1032
rect 33 -1072 45 -1038
rect 413 -1072 425 -1038
rect 33 -1078 425 -1072
rect 491 -1038 883 -1032
rect 491 -1072 503 -1038
rect 871 -1072 883 -1038
rect 491 -1078 883 -1072
<< properties >>
string FIXED_BBOX -1030 -1157 1030 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 2.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
