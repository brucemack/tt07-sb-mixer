magic
tech sky130A
magscale 1 2
timestamp 1715796611
<< metal1 >>
rect 26480 5326 26660 5332
rect 26660 5146 27438 5326
rect 26480 5140 26660 5146
rect 30952 4998 30958 5298
rect 31258 4998 31264 5298
rect 30958 4646 31258 4998
rect 30608 1624 30788 1630
rect 29362 1444 30608 1624
rect 24458 1438 24758 1444
rect 30608 1438 30788 1444
rect 24758 1138 25890 1438
rect 24458 1132 24758 1138
rect 26866 978 27448 1158
rect 26866 760 27046 978
rect 26860 580 26866 760
rect 27046 580 27052 760
<< via1 >>
rect 26480 5146 26660 5326
rect 30958 4998 31258 5298
rect 30608 1444 30788 1624
rect 24458 1138 24758 1438
rect 26866 580 27046 760
<< metal2 >>
rect 30958 5551 31258 5556
rect 26253 5326 26423 5330
rect 26248 5321 26480 5326
rect 26248 5151 26253 5321
rect 26423 5151 26480 5321
rect 26248 5146 26480 5151
rect 26660 5146 26666 5326
rect 30954 5298 30963 5551
rect 31253 5298 31262 5551
rect 30954 5261 30958 5298
rect 31258 5261 31262 5298
rect 26253 5142 26423 5146
rect 30958 4992 31258 4998
rect 30961 1624 31131 1628
rect 30602 1444 30608 1624
rect 30788 1619 31136 1624
rect 30788 1449 30961 1619
rect 31131 1449 31136 1619
rect 30788 1444 31136 1449
rect 24101 1438 24391 1442
rect 30961 1440 31131 1444
rect 24096 1433 24458 1438
rect 24096 1143 24101 1433
rect 24391 1143 24458 1433
rect 24096 1138 24458 1143
rect 24758 1138 24764 1438
rect 24101 1134 24391 1138
rect 26866 760 27046 766
rect 26866 571 27046 580
rect 26862 401 26871 571
rect 27041 401 27050 571
rect 26866 396 27046 401
<< via2 >>
rect 26253 5151 26423 5321
rect 30963 5298 31253 5551
rect 30963 5261 31253 5298
rect 30961 1449 31131 1619
rect 24101 1143 24391 1433
rect 26871 401 27041 571
<< metal3 >>
rect 30958 5861 31258 5862
rect 30953 5563 30959 5861
rect 31257 5563 31263 5861
rect 30958 5551 31258 5563
rect 25901 5326 26079 5331
rect 25900 5325 26428 5326
rect 25900 5147 25901 5325
rect 26079 5321 26428 5325
rect 26079 5151 26253 5321
rect 26423 5151 26428 5321
rect 30958 5261 30963 5551
rect 31253 5261 31258 5551
rect 30958 5256 31258 5261
rect 26079 5147 26428 5151
rect 25900 5146 26428 5147
rect 25901 5141 26079 5146
rect 31283 1624 31461 1629
rect 30956 1623 31462 1624
rect 30956 1619 31283 1623
rect 30956 1449 30961 1619
rect 31131 1449 31283 1619
rect 30956 1445 31283 1449
rect 31461 1445 31462 1623
rect 30956 1444 31462 1445
rect 1645 1438 1943 1443
rect 31283 1439 31461 1444
rect 1644 1437 24396 1438
rect 1644 1139 1645 1437
rect 1943 1433 24396 1437
rect 1943 1143 24101 1433
rect 24391 1143 24396 1433
rect 1943 1139 24396 1143
rect 1644 1138 24396 1139
rect 1645 1133 1943 1138
rect 26866 571 27046 576
rect 26866 401 26871 571
rect 27041 401 27046 571
rect 26866 385 27046 401
rect 26861 207 26867 385
rect 27045 207 27051 385
rect 26866 206 27046 207
<< via3 >>
rect 30959 5563 31257 5861
rect 25901 5147 26079 5325
rect 31283 1445 31461 1623
rect 1645 1139 1943 1437
rect 26867 207 27045 385
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1438 500 44152
rect 9800 6106 10100 44152
rect 9800 5861 31258 6106
rect 9800 5806 30959 5861
rect 200 1437 1944 1438
rect 200 1139 1645 1437
rect 1943 1139 1944 1437
rect 200 1138 1944 1139
rect 200 1000 500 1138
rect 9800 1000 10100 5806
rect 30958 5563 30959 5806
rect 31257 5563 31258 5861
rect 30958 5562 31258 5563
rect 22450 5325 26080 5326
rect 22450 5147 25901 5325
rect 26079 5147 26080 5325
rect 22450 5146 26080 5147
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 5146
rect 31282 1623 31462 1624
rect 31282 1445 31283 1623
rect 31461 1445 31462 1623
rect 26866 385 27046 386
rect 26866 207 26867 385
rect 27045 207 27046 385
rect 26866 0 27046 207
rect 31282 0 31462 1445
use sb_mixer  sb_mixer_0
timestamp 1715793612
transform 0 -1 29296 1 0 446
box 520 -1934 4922 3642
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
