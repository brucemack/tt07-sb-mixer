magic
tech sky130A
magscale 1 2
timestamp 1716640455
<< metal1 >>
rect 20530 8948 20536 9148
rect 20736 8948 20982 9148
rect 20782 7628 20982 8074
rect 26040 7524 26050 7724
rect 26240 7524 26250 7724
rect 20782 7422 20982 7428
rect 26372 4010 26828 4210
rect 27028 4010 27034 4210
rect 31738 2708 31926 2714
rect 31738 2492 31926 2520
rect 30834 2304 31926 2492
rect 24992 1670 25292 1676
rect 25292 1370 25906 1670
rect 24992 1364 25292 1370
<< via1 >>
rect 20536 8948 20736 9148
rect 20782 7428 20982 7628
rect 26050 7524 26240 7724
rect 26828 4010 27028 4210
rect 31738 2520 31926 2708
rect 24992 1370 25292 1670
<< metal2 >>
rect 20536 9148 20736 9154
rect 20293 8948 20302 9148
rect 20502 8948 20536 9148
rect 20536 8942 20736 8948
rect 26050 7724 26240 7734
rect 20782 7628 20982 7637
rect 20776 7428 20782 7628
rect 20982 7428 20988 7628
rect 26050 7514 26240 7524
rect 20782 7419 20982 7428
rect 26828 4210 27028 4216
rect 27028 4010 27062 4210
rect 27262 4010 27271 4210
rect 26828 4004 27028 4010
rect 31738 2910 31926 2919
rect 31738 2708 31926 2722
rect 31732 2520 31738 2708
rect 31926 2520 31932 2708
rect 24681 1670 24971 1674
rect 24676 1665 24992 1670
rect 24676 1375 24681 1665
rect 24971 1375 24992 1665
rect 24676 1370 24992 1375
rect 25292 1370 25298 1670
rect 24681 1366 24971 1370
<< via2 >>
rect 20302 8948 20502 9148
rect 20782 7428 20982 7628
rect 26050 7524 26240 7724
rect 27062 4010 27262 4210
rect 31738 2722 31926 2910
rect 24681 1375 24971 1665
<< metal3 >>
rect 23606 14968 23612 15032
rect 23676 14968 23682 15032
rect 20297 9148 20507 9153
rect 19110 8948 20302 9148
rect 20502 8948 20507 9148
rect 8589 4278 8887 4283
rect 8588 4277 10598 4278
rect 8588 3979 8589 4277
rect 8887 3979 10598 4277
rect 8588 3978 10598 3979
rect 10898 3978 10904 4278
rect 8589 3973 8887 3978
rect 19110 930 19310 8948
rect 20297 8943 20507 8948
rect 23614 7698 23674 14968
rect 26040 7724 26250 7729
rect 26040 7698 26050 7724
rect 23614 7638 26050 7698
rect 20777 7628 20987 7633
rect 20777 7428 20782 7628
rect 20982 7428 20987 7628
rect 26040 7524 26050 7638
rect 26240 7524 26250 7724
rect 26040 7519 26250 7524
rect 20777 7423 20987 7428
rect 20782 7322 20982 7423
rect 20312 7122 20982 7322
rect 20312 1288 20512 7122
rect 27057 4210 27267 4215
rect 27057 4010 27062 4210
rect 27262 4010 31454 4210
rect 27057 4005 27267 4010
rect 24317 1670 24615 1675
rect 24316 1669 24976 1670
rect 24316 1371 24317 1669
rect 24615 1665 24976 1669
rect 24615 1375 24681 1665
rect 24971 1375 24976 1665
rect 24615 1371 24976 1375
rect 24316 1370 24976 1371
rect 24317 1365 24615 1370
rect 20312 1088 27042 1288
rect 19110 730 22660 930
rect 22460 668 22660 730
rect 26842 800 27042 1088
rect 26842 594 27042 600
rect 31254 750 31454 4010
rect 31738 3130 31926 3136
rect 31738 2915 31926 2942
rect 31733 2910 31931 2915
rect 31733 2722 31738 2910
rect 31926 2722 31931 2910
rect 31733 2717 31931 2722
rect 31254 544 31454 550
rect 22460 462 22660 468
<< via3 >>
rect 23612 14968 23676 15032
rect 8589 3979 8887 4277
rect 10598 3978 10898 4278
rect 24317 1371 24615 1669
rect 22460 468 22660 668
rect 26842 600 27042 800
rect 31738 2942 31926 3130
rect 31254 550 31454 750
<< metal4 >>
rect 798 45050 858 45152
rect 796 44952 858 45050
rect 796 44750 856 44952
rect 1534 44750 1594 45152
rect 2270 44750 2330 45152
rect 3006 44750 3066 45152
rect 3742 44750 3802 45152
rect 4478 44750 4538 45152
rect 5214 44750 5274 45152
rect 5950 44750 6010 45152
rect 6686 44750 6746 45152
rect 7422 44750 7482 45152
rect 8158 44750 8218 45152
rect 8894 44750 8954 45152
rect 9630 44750 9690 45152
rect 10366 44750 10426 45152
rect 11102 44750 11162 45152
rect 11838 44750 11898 45152
rect 12574 44750 12634 45152
rect 13310 44750 13370 45152
rect 14046 44750 14106 45152
rect 14782 44750 14842 45152
rect 15518 44750 15578 45152
rect 16254 44750 16314 45152
rect 16990 44750 17050 45152
rect 17726 44750 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 796 44690 17786 44750
rect 1096 44684 1396 44690
rect 3006 44682 3066 44690
rect 3742 44688 4542 44690
rect 5214 44684 5274 44690
rect 5950 44680 6010 44690
rect 8894 44684 8954 44690
rect 200 44110 500 44152
rect 200 43810 504 44110
rect 9046 44022 9106 44690
rect 10366 44684 10426 44690
rect 11102 44688 11162 44690
rect 11838 44688 11898 44690
rect 12574 44678 12634 44690
rect 9800 44022 10100 44152
rect 9046 43962 10100 44022
rect 200 4278 500 43810
rect 9800 14396 10100 43962
rect 23614 15033 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23611 15032 23677 15033
rect 23611 14968 23612 15032
rect 23676 14968 23677 15032
rect 23611 14967 23677 14968
rect 9800 14376 29878 14396
rect 9800 14188 31926 14376
rect 9800 14096 29878 14188
rect 200 4277 8888 4278
rect 200 3979 8589 4277
rect 8887 3979 8888 4277
rect 200 3978 8888 3979
rect 200 1000 500 3978
rect 9800 1000 10100 14096
rect 10597 4278 10899 4279
rect 10597 3978 10598 4278
rect 10898 3978 19002 4278
rect 10597 3977 10899 3978
rect 18702 1670 19002 3978
rect 31738 3131 31926 14188
rect 31737 3130 31927 3131
rect 31737 2942 31738 3130
rect 31926 2942 31927 3130
rect 31737 2941 31927 2942
rect 18702 1669 24616 1670
rect 18702 1371 24317 1669
rect 24615 1371 24616 1669
rect 18702 1370 24616 1371
rect 26841 800 27043 801
rect 22459 668 22661 669
rect 22459 468 22460 668
rect 22660 468 22661 668
rect 26841 600 26842 800
rect 27042 600 27043 800
rect 26841 599 27043 600
rect 31253 750 31455 751
rect 22459 467 22661 468
rect 22460 200 22660 467
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22660 200
rect 22460 -10 22660 0
rect 26842 200 27042 599
rect 31253 550 31254 750
rect 31454 550 31455 750
rect 31253 549 31455 550
rect 31254 200 31454 549
rect 26842 0 27046 200
rect 31254 6 31462 200
rect 31282 0 31462 6
rect 26842 -54 27042 0
use db_mixer  db_mixer_0
timestamp 1716600219
transform 0 -1 26026 1 0 710
box 720 -5014 12418 6460
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
