magic
tech sky130A
magscale 1 2
timestamp 1716650609
<< error_s >>
rect 26230 7668 26300 7748
rect 26200 7662 26300 7668
rect 26048 7616 26300 7662
rect 26048 7606 26248 7616
<< metal1 >>
rect 20530 8948 20536 9148
rect 20736 8948 20982 9148
rect 20782 7628 20982 8074
rect 26038 7606 26048 7662
rect 26248 7606 26258 7662
rect 20782 7422 20982 7428
rect 26372 4010 26828 4210
rect 27028 4010 27034 4210
<< via1 >>
rect 20536 8948 20736 9148
rect 20782 7428 20982 7628
rect 26048 7606 26248 7662
rect 26828 4010 27028 4210
<< metal2 >>
rect 24995 15554 25004 15614
rect 25064 15611 25073 15614
rect 25064 15557 25313 15611
rect 25064 15554 25073 15557
rect 20536 9148 20736 9154
rect 20293 8948 20302 9148
rect 20502 8948 20536 9148
rect 20536 8942 20736 8948
rect 25259 7660 25313 15557
rect 26048 7662 26248 7672
rect 20782 7628 20982 7637
rect 20776 7428 20782 7628
rect 20982 7428 20988 7628
rect 25256 7606 26048 7660
rect 26048 7596 26248 7606
rect 20782 7419 20982 7428
rect 26828 4210 27028 4216
rect 27028 4010 27062 4210
rect 27262 4010 27271 4210
rect 26828 4004 27028 4010
<< via2 >>
rect 25004 15554 25064 15614
rect 20302 8948 20502 9148
rect 20782 7428 20982 7628
rect 27062 4010 27262 4210
<< metal3 >>
rect 23606 41874 23612 41938
rect 23676 41874 23682 41938
rect 23614 41366 23674 41874
rect 23612 41360 23676 41366
rect 23612 41290 23676 41296
rect 23606 16832 23612 16896
rect 23676 16832 23682 16896
rect 23614 16628 23674 16832
rect 23612 16622 23676 16628
rect 23612 16552 23676 16558
rect 24790 15552 24796 15616
rect 24860 15614 24866 15616
rect 24999 15614 25069 15619
rect 24860 15554 25004 15614
rect 25064 15554 25069 15614
rect 24860 15552 24866 15554
rect 24999 15549 25069 15554
rect 20297 9148 20507 9153
rect 19110 8948 20302 9148
rect 20502 8948 20507 9148
rect 8589 4278 8887 4283
rect 8588 4277 10598 4278
rect 8588 3979 8589 4277
rect 8887 3979 10598 4277
rect 8588 3978 10598 3979
rect 10898 3978 10904 4278
rect 8589 3973 8887 3978
rect 19110 930 19310 8948
rect 20297 8943 20507 8948
rect 20777 7628 20987 7633
rect 20777 7428 20782 7628
rect 20982 7428 20987 7628
rect 20777 7423 20987 7428
rect 20782 7322 20982 7423
rect 20312 7122 20982 7322
rect 20312 1288 20512 7122
rect 27057 4210 27267 4215
rect 27057 4010 27062 4210
rect 27262 4010 31454 4210
rect 27057 4005 27267 4010
rect 20312 1088 27042 1288
rect 19110 730 22660 930
rect 22460 668 22660 730
rect 26842 800 27042 1088
rect 26842 594 27042 600
rect 31254 750 31454 4010
rect 31254 544 31454 550
rect 22460 462 22660 468
<< via3 >>
rect 23612 41874 23676 41938
rect 23612 41296 23676 41360
rect 23612 16832 23676 16896
rect 23612 16558 23676 16622
rect 24796 15552 24860 15616
rect 8589 3979 8887 4277
rect 10598 3978 10898 4278
rect 22460 468 22660 668
rect 26842 600 27042 800
rect 31254 550 31454 750
<< metal4 >>
rect 798 45050 858 45152
rect 796 44952 858 45050
rect 796 44750 856 44952
rect 1534 44750 1594 45152
rect 2270 44750 2330 45152
rect 3006 44750 3066 45152
rect 3742 44750 3802 45152
rect 4478 44750 4538 45152
rect 5214 44750 5274 45152
rect 5950 44750 6010 45152
rect 6686 44750 6746 45152
rect 7422 44750 7482 45152
rect 8158 44750 8218 45152
rect 8894 44750 8954 45152
rect 9630 44750 9690 45152
rect 10366 44750 10426 45152
rect 11102 44750 11162 45152
rect 11838 44750 11898 45152
rect 12574 44750 12634 45152
rect 13310 44750 13370 45152
rect 14046 44750 14106 45152
rect 14782 44750 14842 45152
rect 15518 44750 15578 45152
rect 16254 44750 16314 45152
rect 16990 44750 17050 45152
rect 17726 44750 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 796 44690 17786 44750
rect 1096 44684 1396 44690
rect 3006 44682 3066 44690
rect 3742 44688 4542 44690
rect 5214 44684 5274 44690
rect 5950 44680 6010 44690
rect 8894 44684 8954 44690
rect 200 44110 500 44152
rect 200 43810 504 44110
rect 9046 44022 9106 44690
rect 10366 44684 10426 44690
rect 11102 44688 11162 44690
rect 11838 44688 11898 44690
rect 12574 44678 12634 44690
rect 9800 44022 10100 44152
rect 9046 43962 10100 44022
rect 200 4278 500 43810
rect 9800 14396 10100 43962
rect 16990 43638 17050 44690
rect 23614 41939 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23611 41938 23677 41939
rect 23611 41874 23612 41938
rect 23676 41874 23677 41938
rect 23611 41873 23677 41874
rect 23611 41360 23677 41361
rect 23611 41296 23612 41360
rect 23676 41296 23677 41360
rect 23611 41295 23677 41296
rect 23614 16897 23674 41295
rect 23611 16896 23677 16897
rect 23611 16832 23612 16896
rect 23676 16832 23677 16896
rect 23611 16831 23677 16832
rect 23611 16622 23677 16623
rect 23611 16558 23612 16622
rect 23676 16558 23677 16622
rect 23611 16557 23677 16558
rect 23614 15614 23674 16557
rect 24795 15616 24861 15617
rect 24795 15614 24796 15616
rect 23596 15554 24796 15614
rect 23614 15450 23674 15554
rect 24795 15552 24796 15554
rect 24860 15552 24861 15616
rect 24795 15551 24861 15552
rect 9800 14376 29878 14396
rect 9800 14188 29880 14376
rect 9800 14096 29878 14188
rect 200 4277 8888 4278
rect 200 3979 8589 4277
rect 8887 3979 8888 4277
rect 200 3978 8888 3979
rect 200 1000 500 3978
rect 9800 1000 10100 14096
rect 29578 11748 29878 14096
rect 10597 4278 10899 4279
rect 10597 3978 10598 4278
rect 10898 3978 19866 4278
rect 10597 3977 10899 3978
rect 18702 3938 19002 3978
rect 26841 800 27043 801
rect 22459 668 22661 669
rect 22459 468 22460 668
rect 22660 468 22661 668
rect 26841 600 26842 800
rect 27042 600 27043 800
rect 26841 599 27043 600
rect 31253 750 31455 751
rect 22459 467 22661 468
rect 22460 200 22660 467
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22660 200
rect 22460 -10 22660 0
rect 26842 200 27042 599
rect 31253 550 31254 750
rect 31454 550 31455 750
rect 31253 549 31455 550
rect 31254 200 31454 549
rect 26842 0 27046 200
rect 31254 6 31462 200
rect 31282 0 31462 6
rect 26842 -54 27042 0
use db_mixer  db_mixer_0
timestamp 1716650609
transform 0 -1 26026 1 0 710
box 720 -5014 12418 6460
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
