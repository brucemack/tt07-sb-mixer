magic
tech sky130A
magscale 1 2
timestamp 1717070921
<< metal1 >>
rect 20530 8948 20536 9148
rect 20736 8948 20982 9148
rect 20782 7628 20982 8074
rect 20782 7422 20982 7428
rect 26107 7347 26117 7401
rect 26171 7347 26181 7401
rect 26372 4010 26828 4210
rect 27028 4010 27034 4210
<< via1 >>
rect 20536 8948 20736 9148
rect 20782 7428 20982 7628
rect 26117 7347 26171 7401
rect 26828 4010 27028 4210
<< metal2 >>
rect 16990 44256 17050 44258
rect 16983 44200 16992 44256
rect 17048 44200 17057 44256
rect 16990 44108 17050 44200
rect 12850 44048 17050 44108
rect 17726 44078 17786 44080
rect 12850 41464 12910 44048
rect 17719 44022 17728 44078
rect 17784 44022 17793 44078
rect 17726 43886 17786 44022
rect 14778 43826 17786 43886
rect 14778 41356 14838 43826
rect 22878 43822 22938 43824
rect 22871 43766 22880 43822
rect 22936 43766 22945 43822
rect 22878 43564 22938 43766
rect 16720 43504 22938 43564
rect 16720 41536 16780 43504
rect 18644 42404 18704 42406
rect 18637 42348 18646 42404
rect 18702 42348 18711 42404
rect 18644 41534 18704 42348
rect 24995 15554 25004 15614
rect 25064 15611 25073 15614
rect 25064 15557 25313 15611
rect 25064 15554 25073 15557
rect 20536 9148 20736 9154
rect 20293 8948 20302 9148
rect 20502 8948 20536 9148
rect 20536 8942 20736 8948
rect 20782 7628 20982 7637
rect 20776 7428 20782 7628
rect 20982 7428 20988 7628
rect 20782 7419 20982 7428
rect 25259 7401 25313 15557
rect 26117 7401 26171 7411
rect 25259 7347 26117 7401
rect 26117 7337 26171 7347
rect 26828 4210 27028 4216
rect 27028 4010 27062 4210
rect 27262 4010 27271 4210
rect 26828 4004 27028 4010
<< via2 >>
rect 16992 44200 17048 44256
rect 17728 44022 17784 44078
rect 22880 43766 22936 43822
rect 18646 42348 18702 42404
rect 25004 15554 25064 15614
rect 20302 8948 20502 9148
rect 20782 7428 20982 7628
rect 27062 4010 27262 4210
<< metal3 >>
rect 16982 44352 16988 44416
rect 17052 44352 17058 44416
rect 16990 44261 17050 44352
rect 17718 44298 17724 44362
rect 17788 44298 17794 44362
rect 16987 44256 17053 44261
rect 16987 44200 16992 44256
rect 17048 44200 17053 44256
rect 16987 44195 17053 44200
rect 17726 44083 17786 44298
rect 29990 44182 30054 44188
rect 18644 44120 29990 44180
rect 17723 44078 17789 44083
rect 17723 44022 17728 44078
rect 17784 44022 17789 44078
rect 17723 44017 17789 44022
rect 18644 42409 18704 44120
rect 29990 44112 30054 44118
rect 22870 43952 22876 44016
rect 22940 43952 22946 44016
rect 22878 43827 22938 43952
rect 22875 43822 22941 43827
rect 22875 43766 22880 43822
rect 22936 43766 22941 43822
rect 22875 43761 22941 43766
rect 18641 42404 18707 42409
rect 18641 42348 18646 42404
rect 18702 42348 18707 42404
rect 18641 42343 18707 42348
rect 23606 41874 23612 41938
rect 23676 41874 23682 41938
rect 23614 41366 23674 41874
rect 23612 41360 23676 41366
rect 23612 41290 23676 41296
rect 10593 33688 10911 33693
rect 9058 33368 9064 33688
rect 9384 33687 10912 33688
rect 9384 33369 10593 33687
rect 10911 33369 10912 33687
rect 9384 33368 10912 33369
rect 10593 33363 10911 33368
rect 23606 16832 23612 16896
rect 23676 16832 23682 16896
rect 23614 16628 23674 16832
rect 23612 16622 23676 16628
rect 23612 16552 23676 16558
rect 24790 15552 24796 15616
rect 24860 15614 24866 15616
rect 24999 15614 25069 15619
rect 24860 15554 25004 15614
rect 25064 15554 25069 15614
rect 24860 15552 24866 15554
rect 24999 15549 25069 15554
rect 20297 9148 20507 9153
rect 19110 8948 20302 9148
rect 20502 8948 20507 9148
rect 8589 4278 8887 4283
rect 8588 4277 10598 4278
rect 8588 3979 8589 4277
rect 8887 3979 10598 4277
rect 8588 3978 10598 3979
rect 10898 3978 10904 4278
rect 8589 3973 8887 3978
rect 19110 930 19310 8948
rect 20297 8943 20507 8948
rect 20777 7628 20987 7633
rect 20777 7428 20782 7628
rect 20982 7428 20987 7628
rect 20777 7423 20987 7428
rect 20782 7322 20982 7423
rect 20312 7122 20982 7322
rect 20312 1288 20512 7122
rect 27057 4210 27267 4215
rect 27057 4010 27062 4210
rect 27262 4010 31454 4210
rect 27057 4005 27267 4010
rect 20312 1156 27042 1288
rect 20312 1088 27046 1156
rect 19110 730 22660 930
rect 26842 874 27046 1088
rect 22450 688 22660 730
rect 22450 533 22630 688
rect 26866 645 27046 874
rect 31254 750 31454 4010
rect 22445 355 22451 533
rect 22629 355 22635 533
rect 26861 467 26867 645
rect 27045 467 27051 645
rect 31254 544 31454 550
rect 26866 466 27046 467
rect 22450 354 22630 355
<< via3 >>
rect 16988 44352 17052 44416
rect 17724 44298 17788 44362
rect 29990 44118 30054 44182
rect 22876 43952 22940 44016
rect 23612 41874 23676 41938
rect 23612 41296 23676 41360
rect 9064 33368 9384 33688
rect 10593 33369 10911 33687
rect 23612 16832 23676 16896
rect 23612 16558 23676 16622
rect 24796 15552 24860 15616
rect 8589 3979 8887 4277
rect 10598 3978 10898 4278
rect 22451 355 22629 533
rect 26867 467 27045 645
rect 31254 550 31454 750
<< metal4 >>
rect 798 45050 858 45152
rect 796 44952 858 45050
rect 796 44750 856 44952
rect 1534 44750 1594 45152
rect 2270 44750 2330 45152
rect 3006 44750 3066 45152
rect 3742 44750 3802 45152
rect 4478 44750 4538 45152
rect 5214 44750 5274 45152
rect 5950 44750 6010 45152
rect 6686 44750 6746 45152
rect 7422 44750 7482 45152
rect 8158 44750 8218 45152
rect 8894 44750 8954 45152
rect 9630 44750 9690 45152
rect 10366 44750 10426 45152
rect 11102 44750 11162 45152
rect 11838 44750 11898 45152
rect 12574 44750 12634 45152
rect 13310 44750 13370 45152
rect 14046 44750 14106 45152
rect 14782 44750 14842 45152
rect 15518 44750 15578 45152
rect 16254 44750 16314 45152
rect 796 44690 16380 44750
rect 1096 44684 1396 44690
rect 3006 44682 3066 44690
rect 3742 44688 4542 44690
rect 5214 44684 5274 44690
rect 5950 44680 6010 44690
rect 8894 44684 8954 44690
rect 200 44110 500 44152
rect 200 43810 504 44110
rect 9046 44022 9106 44690
rect 10366 44684 10426 44690
rect 11102 44688 11162 44690
rect 11838 44688 11898 44690
rect 12574 44678 12634 44690
rect 16990 44417 17050 45152
rect 16987 44416 17053 44417
rect 16987 44352 16988 44416
rect 17052 44352 17053 44416
rect 17726 44363 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 16987 44351 17053 44352
rect 17723 44362 17789 44363
rect 17723 44298 17724 44362
rect 17788 44298 17789 44362
rect 17723 44297 17789 44298
rect 9800 44022 10100 44152
rect 9046 43962 10100 44022
rect 22878 44017 22938 45152
rect 200 33688 500 43810
rect 9063 33688 9385 33689
rect 180 33368 9064 33688
rect 9384 33368 9385 33688
rect 200 4278 500 33368
rect 9063 33367 9385 33368
rect 9800 32795 10100 43962
rect 22875 44016 22941 44017
rect 22875 43952 22876 44016
rect 22940 43952 22941 44016
rect 22875 43951 22941 43952
rect 23614 41939 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 29989 44182 30055 44183
rect 29989 44118 29990 44182
rect 30054 44180 30055 44182
rect 30238 44180 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 30054 44120 30298 44180
rect 30054 44118 30055 44120
rect 29989 44117 30055 44118
rect 23611 41938 23677 41939
rect 23611 41874 23612 41938
rect 23676 41874 23677 41938
rect 23611 41873 23677 41874
rect 23611 41360 23677 41361
rect 23611 41296 23612 41360
rect 23676 41296 23677 41360
rect 23611 41295 23677 41296
rect 13062 33688 13382 34326
rect 10592 33687 13382 33688
rect 10592 33369 10593 33687
rect 10911 33369 13382 33687
rect 10592 33368 13382 33369
rect 13912 32795 14246 34362
rect 9797 32461 14246 32795
rect 9800 14396 10100 32461
rect 23614 16897 23674 41295
rect 23611 16896 23677 16897
rect 23611 16832 23612 16896
rect 23676 16832 23677 16896
rect 23611 16831 23677 16832
rect 23611 16622 23677 16623
rect 23611 16558 23612 16622
rect 23676 16558 23677 16622
rect 23611 16557 23677 16558
rect 23614 15614 23674 16557
rect 24795 15616 24861 15617
rect 24795 15614 24796 15616
rect 23596 15554 24796 15614
rect 23614 15450 23674 15554
rect 24795 15552 24796 15554
rect 24860 15552 24861 15616
rect 24795 15551 24861 15552
rect 9800 14376 29878 14396
rect 9800 14188 29880 14376
rect 9800 14096 29878 14188
rect 200 4277 8888 4278
rect 200 3979 8589 4277
rect 8887 3979 8888 4277
rect 200 3978 8888 3979
rect 200 1000 500 3978
rect 9800 1000 10100 14096
rect 29578 11748 29878 14096
rect 10597 4278 10899 4279
rect 10597 3978 10598 4278
rect 10898 3978 19866 4278
rect 10597 3977 10899 3978
rect 18702 3938 19002 3978
rect 31253 750 31455 751
rect 26866 645 27046 646
rect 22450 533 22630 534
rect 22450 355 22451 533
rect 22629 355 22630 533
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 355
rect 26866 467 26867 645
rect 27045 467 27046 645
rect 31253 550 31254 750
rect 31454 550 31455 750
rect 31253 549 31455 550
rect 26866 0 27046 467
rect 31254 200 31454 549
rect 31254 6 31462 200
rect 31282 0 31462 6
use db_mixer  db_mixer_0 ~/tt07-sb-mixer/mag
timestamp 1716653920
transform 0 -1 26026 1 0 710
box 720 -5014 12418 6460
use quadrature_divider  quadrature_divider_0
timestamp 1717070208
transform 1 0 11822 0 1 33724
box 514 496 7520 8000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
