magic
tech sky130A
magscale 1 2
timestamp 1715782654
<< pwell >>
rect 3830 1736 4050 1738
rect 3826 1666 4050 1736
rect 3826 1664 4046 1666
<< viali >>
rect 1400 2136 1606 2170
rect 3834 2120 4016 2190
rect 2686 1651 2720 1685
rect 1400 1614 1606 1650
rect 3830 1602 4072 1656
rect 2606 1551 2640 1585
rect 2614 691 2648 725
rect 2694 607 2728 641
rect 1336 272 1682 356
rect 3874 284 4144 350
rect 3756 -1098 3824 -346
<< metal1 >>
rect 776 3630 4002 3642
rect 776 3442 4030 3630
rect 1424 2820 1580 3442
rect 1424 2266 1434 2694
rect 1568 2266 1578 2694
rect 1390 2170 1624 2186
rect 1390 2136 1400 2170
rect 1606 2136 1624 2170
rect 520 1864 1046 2064
rect 1246 1864 1252 2064
rect 1390 1650 1624 2136
rect 2330 2054 2530 2254
rect 1390 1614 1400 1650
rect 1606 1614 1624 1650
rect 1390 1598 1624 1614
rect 2353 1608 2419 2054
rect 2904 1898 3104 3442
rect 3874 2814 4030 3442
rect 2740 1862 3104 1898
rect 2904 1858 3104 1862
rect 3812 2190 4086 2206
rect 3812 2120 3834 2190
rect 4016 2120 4086 2190
rect 2672 1685 2894 1692
rect 2672 1651 2686 1685
rect 2720 1651 2894 1685
rect 2672 1640 2894 1651
rect 2350 1585 2664 1608
rect 1078 1506 2138 1558
rect 2350 1551 2606 1585
rect 2640 1551 2664 1585
rect 2350 1542 2664 1551
rect 2091 1485 2138 1506
rect 2272 1485 2317 1486
rect 2847 1485 2892 1640
rect 1006 486 1016 1474
rect 1072 486 1082 1474
rect 1448 490 1458 1458
rect 1540 490 1550 1458
rect 1922 488 1932 1464
rect 1992 488 2002 1464
rect 2091 1440 2892 1485
rect 2091 446 2138 1440
rect 2186 1302 2784 1368
rect 1080 400 2142 446
rect 1306 356 1720 364
rect 1306 272 1336 356
rect 1682 272 1720 356
rect 1306 235 1720 272
rect 2186 235 2268 1302
rect 2847 1213 2892 1440
rect 2345 1147 2892 1213
rect 2345 742 2411 1147
rect 2976 1052 3048 1858
rect 3812 1656 4086 2120
rect 4254 1864 4260 2064
rect 4460 1864 4922 2064
rect 3812 1602 3830 1656
rect 4072 1602 4086 1656
rect 3812 1582 4086 1602
rect 2550 976 3048 1052
rect 3158 1508 4342 1552
rect 2345 725 2676 742
rect 2345 691 2614 725
rect 2648 691 2676 725
rect 2345 682 2676 691
rect 2345 677 2411 682
rect 3158 654 3218 1508
rect 2678 641 3218 654
rect 2678 607 2694 641
rect 2728 607 3218 641
rect 2678 590 3218 607
rect 2536 235 2812 520
rect 3092 442 3218 590
rect 3420 484 3430 1466
rect 3500 484 3510 1466
rect 3876 488 3886 1466
rect 3974 488 3984 1466
rect 4342 482 4352 1470
rect 4424 482 4434 1470
rect 3092 402 4342 442
rect 3094 398 4342 402
rect 3860 350 4156 356
rect 3860 284 3874 350
rect 4144 284 4156 350
rect 3860 235 4156 284
rect 1302 18 4156 235
rect 1306 14 1720 18
rect 984 -140 1184 -72
rect 974 -182 3618 -140
rect 984 -272 1184 -182
rect 1606 -1262 1634 -182
rect 1802 -1216 1812 -216
rect 1884 -1216 1894 -216
rect 2254 -1206 2264 -222
rect 2344 -1206 2354 -222
rect 2710 -1216 2720 -216
rect 2792 -1216 2802 -216
rect 3164 -1202 3174 -230
rect 3254 -1202 3264 -230
rect 3640 -1200 3650 -218
rect 3706 -1200 3716 -218
rect 3860 -254 4156 18
rect 3744 -346 4156 -254
rect 3744 -1098 3756 -346
rect 3824 -1098 4156 -346
rect 3744 -1150 4156 -1098
rect 1606 -1290 3624 -1262
rect 3902 -1728 4142 -1150
rect 2196 -1928 2202 -1728
rect 2402 -1928 4396 -1728
<< via1 >>
rect 1434 2266 1568 2694
rect 1046 1864 1246 2064
rect 1016 486 1072 1474
rect 1458 490 1540 1458
rect 1932 488 1992 1464
rect 4260 1864 4460 2064
rect 3430 484 3500 1466
rect 3886 488 3974 1466
rect 4352 482 4424 1470
rect 1812 -1216 1884 -216
rect 2264 -1206 2344 -222
rect 2720 -1216 2792 -216
rect 3174 -1202 3254 -230
rect 3650 -1200 3706 -218
rect 2202 -1928 2402 -1728
<< metal2 >>
rect 1434 2694 1568 2704
rect 1568 2266 1570 2286
rect 1046 2064 1246 2070
rect 1434 2064 1570 2266
rect 1246 1864 1570 2064
rect 1046 1858 1246 1864
rect 1434 1722 1570 1864
rect 3856 2064 3998 2690
rect 4260 2064 4460 2070
rect 3856 1864 4260 2064
rect 1016 1474 1072 1484
rect 1462 1468 1542 1722
rect 3856 1716 3998 1864
rect 4260 1858 4460 1864
rect 3898 1476 3954 1716
rect 1016 476 1072 486
rect 1458 1458 1542 1468
rect 1540 1456 1542 1458
rect 1932 1464 1992 1474
rect 1458 480 1540 490
rect 1932 478 1992 488
rect 3430 1466 3500 1476
rect 1022 190 1062 476
rect 1944 190 1984 478
rect 3430 474 3500 484
rect 3886 1466 3974 1476
rect 3886 478 3974 488
rect 4352 1470 4424 1480
rect 4424 482 4426 496
rect 3436 190 3498 474
rect 4352 472 4426 482
rect 4364 190 4426 472
rect 1022 134 4426 190
rect 1026 128 4426 134
rect 1026 88 4424 128
rect 1808 -206 1864 88
rect 2722 -206 2778 88
rect 1808 -216 1884 -206
rect 1808 -288 1812 -216
rect 2264 -222 2344 -212
rect 2264 -1216 2344 -1206
rect 2720 -216 2792 -206
rect 3656 -208 3712 88
rect 3650 -218 3712 -208
rect 3174 -230 3254 -220
rect 3174 -1212 3254 -1202
rect 3706 -288 3712 -218
rect 3650 -1210 3706 -1200
rect 1812 -1226 1884 -1216
rect 2276 -1504 2330 -1216
rect 2720 -1226 2792 -1216
rect 2202 -1522 2402 -1504
rect 3182 -1522 3236 -1212
rect 2202 -1576 3236 -1522
rect 2202 -1728 2402 -1576
rect 2202 -1934 2402 -1928
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2526 0 1 1336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1704896540
transform 1 0 2534 0 1 476
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_lvt_WWWVRA  XM1
timestamp 1715647744
transform 1 0 2759 0 1 -714
box -1083 -710 1083 710
use sky130_fd_pr__nfet_01v8_L3FTKF  XM2
timestamp 1715647744
transform 1 0 1503 0 1 976
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_L3FTKF  XM3
timestamp 1715647744
transform 1 0 3929 0 1 976
box -625 -710 625 710
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR1
timestamp 1715647744
transform 1 0 1503 0 1 2751
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR2
timestamp 1715647744
transform 1 0 3929 0 1 2751
box -235 -651 235 651
<< labels >>
flabel metal1 520 1864 720 2064 0 FreeSans 256 0 0 0 IFOUT_P
port 0 nsew
flabel metal1 4722 1864 4922 2064 0 FreeSans 256 0 0 0 IFOUT_N
port 1 nsew
flabel metal1 984 -272 1184 -72 0 FreeSans 256 0 0 0 RFIN
port 2 nsew
flabel metal1 776 3442 976 3642 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 4196 -1928 4396 -1728 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 2330 2054 2530 2254 0 FreeSans 256 0 0 0 LOIN
port 5 nsew
flabel metal2 1026 88 4424 190 0 FreeSans 1600 0 0 0 v1
flabel metal2 1026 88 4424 190 0 FreeSans 1600 0 0 0 V1
<< end >>
