magic
tech sky130A
magscale 1 2
timestamp 1716495612
<< pwell >>
rect -1083 -710 1083 710
<< nmos >>
rect -887 -500 -487 500
rect -429 -500 -29 500
rect 29 -500 429 500
rect 487 -500 887 500
<< ndiff >>
rect -945 488 -887 500
rect -945 -488 -933 488
rect -899 -488 -887 488
rect -945 -500 -887 -488
rect -487 488 -429 500
rect -487 -488 -475 488
rect -441 -488 -429 488
rect -487 -500 -429 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 429 488 487 500
rect 429 -488 441 488
rect 475 -488 487 488
rect 429 -500 487 -488
rect 887 488 945 500
rect 887 -488 899 488
rect 933 -488 945 488
rect 887 -500 945 -488
<< ndiffc >>
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
<< psubdiff >>
rect -1047 640 -951 674
rect 951 640 1047 674
rect -1047 578 -1013 640
rect 1013 578 1047 640
rect -1047 -640 -1013 -578
rect 1013 -640 1047 -578
rect -1047 -674 -951 -640
rect 951 -674 1047 -640
<< psubdiffcont >>
rect -951 640 951 674
rect -1047 -578 -1013 578
rect 1013 -578 1047 578
rect -951 -674 951 -640
<< poly >>
rect -887 572 -487 588
rect -887 538 -871 572
rect -503 538 -487 572
rect -887 500 -487 538
rect -429 572 -29 588
rect -429 538 -413 572
rect -45 538 -29 572
rect -429 500 -29 538
rect 29 572 429 588
rect 29 538 45 572
rect 413 538 429 572
rect 29 500 429 538
rect 487 572 887 588
rect 487 538 503 572
rect 871 538 887 572
rect 487 500 887 538
rect -887 -538 -487 -500
rect -887 -572 -871 -538
rect -503 -572 -487 -538
rect -887 -588 -487 -572
rect -429 -538 -29 -500
rect -429 -572 -413 -538
rect -45 -572 -29 -538
rect -429 -588 -29 -572
rect 29 -538 429 -500
rect 29 -572 45 -538
rect 413 -572 429 -538
rect 29 -588 429 -572
rect 487 -538 887 -500
rect 487 -572 503 -538
rect 871 -572 887 -538
rect 487 -588 887 -572
<< polycont >>
rect -871 538 -503 572
rect -413 538 -45 572
rect 45 538 413 572
rect 503 538 871 572
rect -871 -572 -503 -538
rect -413 -572 -45 -538
rect 45 -572 413 -538
rect 503 -572 871 -538
<< locali >>
rect -1047 640 -951 674
rect 951 640 1047 674
rect -1047 578 -1013 640
rect 1013 578 1047 640
rect -887 538 -871 572
rect -503 538 -487 572
rect -429 538 -413 572
rect -45 538 -29 572
rect 29 538 45 572
rect 413 538 429 572
rect 487 538 503 572
rect 871 538 887 572
rect -933 488 -899 504
rect -933 -504 -899 -488
rect -475 488 -441 504
rect -475 -504 -441 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 441 488 475 504
rect 441 -504 475 -488
rect 899 488 933 504
rect 899 -504 933 -488
rect -887 -572 -871 -538
rect -503 -572 -487 -538
rect -429 -572 -413 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 413 -572 429 -538
rect 487 -572 503 -538
rect 871 -572 887 -538
rect -1047 -640 -1013 -578
rect 1013 -640 1047 -578
rect -1047 -674 -951 -640
rect 951 -674 1047 -640
<< viali >>
rect -871 538 -503 572
rect -413 538 -45 572
rect 45 538 413 572
rect 503 538 871 572
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
rect -871 -572 -503 -538
rect -413 -572 -45 -538
rect 45 -572 413 -538
rect 503 -572 871 -538
<< metal1 >>
rect -883 572 -491 578
rect -883 538 -871 572
rect -503 538 -491 572
rect -883 532 -491 538
rect -425 572 -33 578
rect -425 538 -413 572
rect -45 538 -33 572
rect -425 532 -33 538
rect 33 572 425 578
rect 33 538 45 572
rect 413 538 425 572
rect 33 532 425 538
rect 491 572 883 578
rect 491 538 503 572
rect 871 538 883 572
rect 491 532 883 538
rect -939 488 -893 500
rect -939 -488 -933 488
rect -899 -488 -893 488
rect -939 -500 -893 -488
rect -481 488 -435 500
rect -481 -488 -475 488
rect -441 -488 -435 488
rect -481 -500 -435 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 435 488 481 500
rect 435 -488 441 488
rect 475 -488 481 488
rect 435 -500 481 -488
rect 893 488 939 500
rect 893 -488 899 488
rect 933 -488 939 488
rect 893 -500 939 -488
rect -883 -538 -491 -532
rect -883 -572 -871 -538
rect -503 -572 -491 -538
rect -883 -578 -491 -572
rect -425 -538 -33 -532
rect -425 -572 -413 -538
rect -45 -572 -33 -538
rect -425 -578 -33 -572
rect 33 -538 425 -532
rect 33 -572 45 -538
rect 413 -572 425 -538
rect 33 -578 425 -572
rect 491 -538 883 -532
rect 491 -572 503 -538
rect 871 -572 883 -538
rect 491 -578 883 -572
<< properties >>
string FIXED_BBOX -1030 -657 1030 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 2.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
