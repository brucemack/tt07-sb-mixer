magic
tech sky130A
magscale 1 2
timestamp 1716650609
<< pwell >>
rect 3478 -550 3886 -394
rect 2700 -2286 2824 -944
rect 2174 -2664 3870 -2522
rect 2174 -2814 3536 -2664
rect 2174 -2848 2308 -2814
rect 3214 -2816 3536 -2814
rect 2172 -3008 2308 -2970
rect 3372 -3008 3534 -2970
rect 2172 -3270 3534 -3008
rect 2172 -3300 2276 -3270
rect 3234 -3300 3534 -3270
rect 2172 -3450 2282 -3420
rect 2172 -3458 3230 -3450
rect 2172 -3720 3532 -3458
rect 2172 -3756 2304 -3720
rect 2172 -3916 2304 -3878
rect 3216 -3916 3530 -3878
rect 2172 -4178 3530 -3916
rect 6314 -4036 8702 -3786
rect 6314 -4100 6672 -4036
rect 8572 -4100 8702 -4036
rect 2172 -4220 2264 -4178
rect 3248 -4220 3530 -4178
rect 6316 -4318 6672 -4248
rect 8572 -4318 8704 -4248
rect 6316 -4562 8704 -4318
<< ndiff >>
rect 3042 -3346 3100 -3334
<< viali >>
rect 5598 4984 5678 5244
rect 9802 5062 9872 5282
rect 4698 3770 5170 3836
rect 6478 3776 6976 3846
rect 8266 3770 8762 3848
rect 10234 3788 10740 3868
rect 12014 3604 12106 3744
rect 2868 3058 2952 3300
rect 7642 31 7676 65
rect 7562 -137 7596 -103
rect 6032 -598 6108 -162
rect 6916 -260 7028 -216
rect 9138 -594 9202 -194
rect 7642 -1169 7676 -1135
rect 7562 -1337 7596 -1303
rect 2270 -4442 2964 -4362
rect 12140 -4426 12300 -4346
rect 7374 -4782 7682 -4706
<< metal1 >>
rect 9562 6398 9756 6400
rect 5714 6370 5936 6378
rect 5714 6198 5736 6370
rect 5930 6198 5940 6370
rect 9548 6202 9558 6398
rect 9754 6202 9764 6398
rect 5714 5558 5936 6198
rect 9562 5494 9756 6202
rect 5394 5244 5696 5260
rect 5394 5190 5598 5244
rect 5312 5020 5322 5190
rect 5494 5020 5598 5190
rect 5394 4984 5598 5020
rect 5678 4984 5696 5244
rect 5394 4972 5696 4984
rect 5724 4622 5914 5398
rect 7164 4622 7364 5244
rect 4042 4426 7754 4622
rect 2584 3716 2594 3908
rect 2922 3716 2932 3908
rect 2704 3028 2808 3716
rect 4042 3610 4238 4426
rect 5724 4424 5914 4426
rect 7212 4292 7420 4298
rect 4834 3900 4844 4082
rect 4686 3874 4844 3900
rect 5018 3900 5028 4082
rect 6628 3902 6638 4084
rect 5018 3874 5184 3900
rect 4686 3836 5184 3874
rect 4686 3770 4698 3836
rect 5170 3770 5184 3836
rect 4686 3760 5184 3770
rect 6460 3866 6638 3902
rect 6830 3902 6840 4084
rect 6830 3866 6988 3902
rect 6460 3846 6988 3866
rect 6460 3776 6478 3846
rect 6976 3776 6988 3846
rect 6460 3756 6988 3776
rect 4452 3610 4758 3620
rect 6892 3614 7176 3618
rect 7212 3614 7420 4084
rect 4042 3414 4758 3610
rect 2856 3300 3106 3308
rect 2856 3058 2868 3300
rect 2952 3294 3106 3300
rect 2952 3086 2994 3294
rect 3168 3086 3178 3294
rect 2952 3058 3106 3086
rect 2856 3022 3106 3058
rect 4452 1678 4758 3414
rect 5108 1870 5428 3614
rect 6230 1870 6560 3610
rect 5108 1680 6560 1870
rect 5356 1674 6560 1680
rect 6892 3406 7420 3614
rect 7558 3600 7754 4426
rect 7858 4292 8066 4298
rect 8238 4292 8438 5244
rect 9546 4456 9750 5402
rect 9790 5282 9994 5294
rect 9790 5062 9802 5282
rect 9872 5188 9994 5282
rect 9872 5106 9944 5188
rect 10040 5106 10050 5188
rect 9872 5062 9994 5106
rect 9790 5044 9994 5062
rect 9544 4292 9752 4456
rect 8066 4285 9752 4292
rect 8066 4099 11407 4285
rect 8066 4084 9752 4099
rect 7858 4078 8066 4084
rect 8406 3912 8416 4056
rect 8254 3878 8416 3912
rect 8610 3912 8620 4056
rect 10328 3912 10338 4046
rect 8610 3878 8774 3912
rect 8254 3848 8774 3878
rect 8254 3770 8266 3848
rect 8762 3770 8774 3848
rect 10218 3898 10338 3912
rect 10586 3912 10596 4046
rect 10586 3898 10752 3912
rect 10218 3868 10752 3898
rect 10218 3788 10234 3868
rect 10740 3788 10752 3868
rect 10218 3776 10752 3788
rect 8254 3756 8774 3770
rect 8028 3600 8356 3630
rect 4756 1406 5106 1632
rect 4756 1056 5165 1406
rect 5515 1056 5521 1406
rect 720 110 908 310
rect 1108 110 1114 310
rect 5694 48 5886 1674
rect 6892 1664 7176 3406
rect 7558 3404 8356 3600
rect 8028 1672 8356 3404
rect 8696 1884 8976 3618
rect 10022 1884 10296 3630
rect 8696 1722 10296 1884
rect 8696 1684 8976 1722
rect 6550 1240 6890 1624
rect 8344 1240 8682 1624
rect 6548 1088 8688 1240
rect 6033 269 6039 619
rect 6389 414 6855 619
rect 6389 298 7940 414
rect 6389 269 6855 298
rect 7122 224 7554 236
rect 7112 136 7122 224
rect 7248 136 7554 224
rect 7842 76 7940 298
rect 3924 -210 5886 48
rect 7630 65 7944 76
rect 7630 31 7642 65
rect 7676 31 7944 65
rect 7630 20 7944 31
rect 6536 -58 6736 -16
rect 6536 -78 7022 -58
rect 6536 -103 7626 -78
rect 6536 -137 7562 -103
rect 7596 -137 7626 -103
rect 6536 -146 7626 -137
rect 6018 -162 6324 -146
rect 3300 -394 3500 -346
rect 3826 -394 5988 -238
rect 3300 -546 5988 -394
rect 3478 -550 5988 -546
rect 3826 -578 5988 -550
rect 6018 -598 6032 -162
rect 6108 -286 6324 -162
rect 6536 -174 7022 -146
rect 6536 -182 6826 -174
rect 6536 -216 6736 -182
rect 6896 -274 6906 -204
rect 7038 -274 7048 -204
rect 6108 -470 6254 -286
rect 6412 -470 6422 -286
rect 7144 -398 7154 -302
rect 7254 -304 7264 -302
rect 7254 -398 7666 -304
rect 7154 -400 7666 -398
rect 6108 -598 6324 -470
rect 7876 -572 7932 20
rect 3932 -828 5886 -606
rect 6018 -610 6324 -598
rect 7110 -628 7932 -572
rect 2700 -1805 2824 -944
rect 2700 -1947 3867 -1805
rect 2700 -2244 2824 -1947
rect 2284 -2484 3224 -2244
rect 3725 -2522 3867 -1947
rect 5680 -1900 5878 -828
rect 7110 -1290 7166 -628
rect 7312 -1056 7934 -962
rect 8062 -1056 8072 -962
rect 8306 -1050 8474 1088
rect 9346 32 9638 1722
rect 10022 1706 10296 1722
rect 10668 3588 10942 3628
rect 11221 3588 11407 4099
rect 12038 4018 12048 4172
rect 12382 4018 12392 4172
rect 11916 3744 12118 3752
rect 11916 3724 12014 3744
rect 11832 3634 11842 3724
rect 11952 3634 12014 3724
rect 11916 3604 12014 3634
rect 12106 3604 12118 3744
rect 10668 3402 11412 3588
rect 11916 3586 12118 3604
rect 10668 1700 10942 3402
rect 12156 3266 12270 4018
rect 9723 1406 10073 1412
rect 10316 1406 10638 1630
rect 10073 1056 10638 1406
rect 9723 1050 10073 1056
rect 10316 1054 10638 1056
rect 9346 -106 11304 32
rect 8986 -194 9210 -182
rect 8986 -296 9138 -194
rect 8844 -496 8854 -296
rect 9066 -496 9138 -296
rect 8986 -594 9138 -496
rect 9202 -594 9210 -194
rect 9356 -204 11304 -106
rect 9246 -238 11408 -232
rect 12150 -238 12300 1294
rect 9246 -552 12300 -238
rect 9246 -564 11408 -552
rect 8986 -612 9210 -594
rect 9360 -822 11298 -592
rect 8306 -1118 8468 -1050
rect 7632 -1135 8468 -1118
rect 7632 -1169 7642 -1135
rect 7676 -1169 8468 -1135
rect 7632 -1184 8468 -1169
rect 8306 -1186 8468 -1184
rect 7110 -1303 7610 -1290
rect 7110 -1337 7562 -1303
rect 7596 -1337 7610 -1303
rect 7110 -1346 7610 -1337
rect 7126 -1600 7136 -1506
rect 7242 -1600 7666 -1506
rect 7138 -1602 7666 -1600
rect 9403 -1900 9601 -822
rect 12150 -1894 12300 -552
rect 5680 -2098 9601 -1900
rect 2174 -2664 3870 -2522
rect 7467 -2564 7665 -2098
rect 2174 -2814 3536 -2664
rect 2174 -2848 2308 -2814
rect 3214 -2816 3536 -2814
rect 2366 -2856 3152 -2852
rect 2366 -2952 2654 -2856
rect 2860 -2952 3152 -2856
rect 2366 -2958 3152 -2952
rect 2172 -3008 2308 -2970
rect 3372 -2999 3534 -2970
rect 3725 -2999 3867 -2664
rect 6656 -2838 8598 -2564
rect 6314 -2981 8702 -2874
rect 3372 -3008 3867 -2999
rect 2172 -3141 3867 -3008
rect 2172 -3270 3534 -3141
rect 2172 -3300 2276 -3270
rect 3234 -3300 3534 -3270
rect 3725 -3304 3867 -3141
rect 5951 -3123 8702 -2981
rect 2322 -3338 2996 -3308
rect 2290 -3388 2996 -3338
rect 2322 -3394 2996 -3388
rect 3140 -3338 3200 -3308
rect 3140 -3388 3234 -3338
rect 3140 -3394 3200 -3388
rect 2322 -3396 3200 -3394
rect 3716 -3404 3726 -3304
rect 3862 -3404 3872 -3304
rect 2172 -3450 2282 -3420
rect 2172 -3458 3230 -3450
rect 2172 -3459 3532 -3458
rect 3725 -3459 3867 -3404
rect 2172 -3601 3867 -3459
rect 2172 -3720 3532 -3601
rect 2172 -3756 2304 -3720
rect 2648 -3768 2658 -3764
rect 2372 -3872 2658 -3768
rect 2864 -3768 2874 -3764
rect 2864 -3872 3152 -3768
rect 2172 -3916 2304 -3878
rect 2372 -3882 3152 -3872
rect 3216 -3916 3530 -3878
rect 2172 -4035 3530 -3916
rect 3725 -4035 3867 -3601
rect 5951 -3415 6093 -3123
rect 6314 -3148 8702 -3123
rect 6314 -3188 6672 -3148
rect 8564 -3188 8702 -3148
rect 7366 -3198 7376 -3194
rect 6740 -3322 7376 -3198
rect 7680 -3198 7690 -3194
rect 7680 -3322 8534 -3198
rect 6314 -3386 6672 -3330
rect 8564 -3386 8702 -3330
rect 6314 -3415 8702 -3386
rect 5951 -3557 8702 -3415
rect 9032 -3476 9128 -2098
rect 5951 -3859 6093 -3557
rect 6314 -3586 8702 -3557
rect 9026 -3572 9032 -3476
rect 9128 -3572 9134 -3476
rect 6314 -3644 6656 -3586
rect 8574 -3644 8702 -3586
rect 6730 -3662 8532 -3660
rect 6730 -3776 7880 -3662
rect 7870 -3778 7880 -3776
rect 8230 -3776 8532 -3662
rect 8230 -3778 8240 -3776
rect 6314 -3832 6656 -3786
rect 8574 -3832 8702 -3786
rect 6314 -3859 8702 -3832
rect 5951 -4001 8702 -3859
rect 12152 -3910 12286 -3832
rect 5951 -4035 6093 -4001
rect 2172 -4078 6093 -4035
rect 2172 -4177 3762 -4078
rect 2172 -4178 3530 -4177
rect 3756 -4178 3762 -4177
rect 3862 -4177 6093 -4078
rect 6314 -4036 8702 -4001
rect 6314 -4100 6672 -4036
rect 8572 -4100 8702 -4036
rect 7362 -4112 7372 -4104
rect 3862 -4178 3868 -4177
rect 2172 -4220 2264 -4178
rect 3248 -4220 3530 -4178
rect 2304 -4320 2988 -4232
rect 3116 -4320 3212 -4232
rect 5951 -4333 6093 -4177
rect 6744 -4236 7372 -4112
rect 7684 -4112 7694 -4104
rect 7684 -4236 8514 -4112
rect 12142 -4174 12152 -3910
rect 12286 -4174 12296 -3910
rect 6744 -4244 8514 -4236
rect 6316 -4318 6672 -4248
rect 8572 -4318 8704 -4248
rect 12152 -4300 12286 -4174
rect 6316 -4333 8704 -4318
rect 2260 -4352 2976 -4348
rect 2260 -4362 2550 -4352
rect 2692 -4362 2976 -4352
rect 2260 -4442 2270 -4362
rect 2964 -4442 2976 -4362
rect 2260 -4456 2550 -4442
rect 2692 -4456 2976 -4442
rect 2260 -4470 2976 -4456
rect 5951 -4475 8704 -4333
rect 12124 -4336 12322 -4328
rect 12124 -4346 12156 -4336
rect 12286 -4346 12322 -4336
rect 12124 -4426 12140 -4346
rect 12300 -4426 12322 -4346
rect 12124 -4452 12156 -4426
rect 12286 -4452 12322 -4426
rect 12124 -4470 12322 -4452
rect 6316 -4522 8704 -4475
rect 6316 -4562 6660 -4522
rect 8570 -4562 8704 -4522
rect 6746 -4580 8524 -4576
rect 6746 -4670 7888 -4580
rect 8246 -4670 8524 -4580
rect 1594 -5008 1782 -4808
rect 1982 -5008 1988 -4808
rect 7344 -4824 7354 -4698
rect 7706 -4824 7716 -4698
<< via1 >>
rect 5736 6198 5930 6370
rect 9558 6202 9754 6398
rect 5322 5020 5494 5190
rect 2594 3716 2922 3908
rect 7212 4084 7420 4292
rect 4844 3874 5018 4082
rect 6638 3866 6830 4084
rect 2994 3086 3168 3294
rect 9944 5106 10040 5188
rect 7858 4084 8066 4292
rect 8416 3878 8610 4056
rect 10338 3898 10586 4046
rect 5165 1056 5515 1406
rect 908 110 1108 310
rect 6039 269 6389 619
rect 7122 136 7248 224
rect 6906 -216 7038 -204
rect 6906 -260 6916 -216
rect 6916 -260 7028 -216
rect 7028 -260 7038 -216
rect 6906 -274 7038 -260
rect 6254 -470 6412 -286
rect 7154 -398 7254 -302
rect 7934 -1056 8062 -962
rect 12048 4018 12382 4172
rect 11842 3634 11952 3724
rect 9723 1056 10073 1406
rect 8854 -496 9066 -296
rect 7136 -1600 7242 -1506
rect 2654 -2952 2860 -2856
rect 2996 -3394 3140 -3308
rect 3726 -3404 3862 -3304
rect 2658 -3872 2864 -3764
rect 7376 -3322 7680 -3194
rect 9032 -3572 9128 -3476
rect 7880 -3778 8230 -3662
rect 3762 -4178 3862 -4078
rect 2988 -4320 3116 -4232
rect 7372 -4236 7684 -4104
rect 12152 -4174 12286 -3910
rect 2550 -4362 2692 -4352
rect 2550 -4442 2692 -4362
rect 2550 -4456 2692 -4442
rect 12156 -4346 12286 -4336
rect 12156 -4426 12286 -4346
rect 12156 -4452 12286 -4426
rect 7888 -4670 8246 -4580
rect 1782 -5008 1982 -4808
rect 7354 -4706 7706 -4698
rect 7354 -4782 7374 -4706
rect 7374 -4782 7682 -4706
rect 7682 -4782 7706 -4706
rect 7354 -4824 7706 -4782
<< metal2 >>
rect 9558 6398 9754 6408
rect 5736 6370 5930 6380
rect 5736 6188 5930 6198
rect 9558 6192 9754 6202
rect 5322 5190 5494 5200
rect 9944 5188 10040 5198
rect 9944 5096 10040 5106
rect 5322 5010 5494 5020
rect 4844 4082 5018 4092
rect 2594 3908 2922 3918
rect 4844 3864 5018 3874
rect 6638 4084 6830 4094
rect 7206 4084 7212 4292
rect 7420 4084 7858 4292
rect 8066 4084 8072 4292
rect 12048 4172 12382 4182
rect 8416 4056 8610 4066
rect 10338 4046 10586 4056
rect 12048 4008 12382 4018
rect 10338 3888 10586 3898
rect 8416 3868 8610 3878
rect 6638 3856 6830 3866
rect 2594 3706 2922 3716
rect 11842 3724 11952 3734
rect 11842 3624 11952 3634
rect 2994 3294 3168 3304
rect 2994 3076 3168 3086
rect 5165 1406 5515 1412
rect 5515 1056 9723 1406
rect 10073 1056 10079 1406
rect 5165 1050 5515 1056
rect 6039 619 6389 1056
rect 908 310 1108 316
rect 1276 110 1285 310
rect 6039 263 6389 269
rect 7122 224 7248 234
rect 7122 126 7248 136
rect 908 104 1108 110
rect 6906 -204 7038 -194
rect 6254 -286 6412 -276
rect 6906 -284 7038 -274
rect 7154 -302 7254 -292
rect 7154 -408 7254 -398
rect 8854 -296 9066 -286
rect 6254 -480 6412 -470
rect 8854 -506 9066 -496
rect 7934 -962 8062 -952
rect 7934 -1066 8062 -1056
rect 7136 -1506 7242 -1496
rect 7136 -1610 7242 -1600
rect 2654 -2856 2860 -2846
rect 2654 -2962 2860 -2952
rect 7376 -3194 7680 -3184
rect 2996 -3302 3140 -3298
rect 3726 -3302 3862 -3294
rect 2996 -3304 3870 -3302
rect 2996 -3308 3726 -3304
rect 3140 -3394 3726 -3308
rect 2996 -3404 3726 -3394
rect 3862 -3404 3870 -3304
rect 7376 -3332 7680 -3322
rect 3726 -3414 3862 -3404
rect 9032 -3476 9128 -3470
rect 7880 -3662 8230 -3652
rect 9032 -3662 9128 -3572
rect 2658 -3764 2864 -3754
rect 8230 -3778 9136 -3662
rect 7880 -3788 9136 -3778
rect 7882 -3792 9136 -3788
rect 2658 -3882 2864 -3872
rect 3762 -4078 3862 -4072
rect 2988 -4228 3116 -4222
rect 3762 -4228 3862 -4178
rect 2988 -4232 3862 -4228
rect 3116 -4320 3862 -4232
rect 7372 -4104 7684 -4094
rect 7372 -4246 7684 -4236
rect 2988 -4328 3862 -4320
rect 2988 -4330 3116 -4328
rect 2550 -4352 2692 -4342
rect 2550 -4466 2692 -4456
rect 7888 -4580 8246 -4570
rect 9032 -4582 9128 -3792
rect 12152 -3910 12286 -3900
rect 12152 -4184 12286 -4174
rect 12156 -4336 12286 -4326
rect 12156 -4462 12286 -4452
rect 8246 -4670 9136 -4582
rect 7888 -4678 9136 -4670
rect 7354 -4688 7706 -4678
rect 7888 -4680 8246 -4678
rect 1782 -4808 1982 -4802
rect 1982 -5008 2002 -4808
rect 2202 -5008 2211 -4808
rect 7354 -4834 7706 -4824
rect 1782 -5014 1982 -5008
<< via2 >>
rect 5736 6198 5930 6370
rect 9558 6202 9754 6398
rect 5322 5020 5494 5190
rect 9944 5106 10040 5188
rect 2594 3716 2922 3908
rect 4844 3874 5018 4082
rect 6638 3866 6830 4084
rect 8416 3878 8610 4056
rect 10338 3898 10586 4046
rect 12048 4018 12382 4172
rect 11842 3634 11952 3724
rect 2994 3086 3168 3294
rect 1076 110 1108 310
rect 1108 110 1276 310
rect 7122 136 7248 224
rect 6906 -274 7038 -204
rect 6254 -470 6412 -286
rect 7154 -398 7254 -302
rect 8854 -496 9066 -296
rect 7934 -1056 8062 -962
rect 7136 -1600 7242 -1506
rect 2654 -2952 2860 -2856
rect 7376 -3322 7680 -3194
rect 2658 -3872 2864 -3764
rect 7372 -4236 7684 -4104
rect 2550 -4456 2692 -4352
rect 12152 -4174 12286 -3910
rect 12156 -4452 12286 -4336
rect 7354 -4698 7706 -4688
rect 2002 -5008 2202 -4808
rect 7354 -4824 7706 -4698
<< metal3 >>
rect 9548 6398 9764 6403
rect 5726 6370 5940 6375
rect 5726 6198 5736 6370
rect 5930 6198 5940 6370
rect 5726 6193 5940 6198
rect 9548 6202 9558 6398
rect 9754 6202 9764 6398
rect 9548 6197 9764 6202
rect 5312 5190 5504 5195
rect 5312 5020 5322 5190
rect 5494 5020 5504 5190
rect 9934 5188 10050 5193
rect 9934 5106 9944 5188
rect 10040 5106 10050 5188
rect 9934 5101 10050 5106
rect 5312 5015 5504 5020
rect 12038 4172 12392 4177
rect 4834 4082 5028 4087
rect 2584 3908 2932 3913
rect 2584 3716 2594 3908
rect 2922 3716 2932 3908
rect 4834 3874 4844 4082
rect 5018 3874 5028 4082
rect 4834 3869 5028 3874
rect 6628 4084 6840 4089
rect 6628 3866 6638 4084
rect 6830 3866 6840 4084
rect 8406 4056 8620 4061
rect 8406 3878 8416 4056
rect 8610 3878 8620 4056
rect 10328 4046 10596 4051
rect 10328 3898 10338 4046
rect 10586 3898 10596 4046
rect 12038 4018 12048 4172
rect 12382 4018 12392 4172
rect 12038 4013 12392 4018
rect 10328 3893 10596 3898
rect 8406 3873 8620 3878
rect 6628 3861 6840 3866
rect 2584 3711 2932 3716
rect 11832 3724 11962 3729
rect 11832 3634 11842 3724
rect 11952 3634 11962 3724
rect 11832 3629 11962 3634
rect 2984 3294 3178 3299
rect 2984 3086 2994 3294
rect 3168 3086 3178 3294
rect 2984 3081 3178 3086
rect 1071 310 1281 315
rect 1071 110 1076 310
rect 1446 110 1452 310
rect 7112 224 7258 229
rect 7112 136 7122 224
rect 7248 136 7258 224
rect 7112 131 7258 136
rect 1071 105 1281 110
rect 6896 -204 7048 -199
rect 6896 -274 6906 -204
rect 7038 -274 7048 -204
rect 6896 -279 7048 -274
rect 6244 -286 6422 -281
rect 6244 -470 6254 -286
rect 6412 -470 6422 -286
rect 8844 -296 9076 -291
rect 7144 -302 7264 -297
rect 7144 -398 7154 -302
rect 7254 -398 7264 -302
rect 7144 -403 7264 -398
rect 6244 -475 6422 -470
rect 8844 -496 8854 -296
rect 9066 -496 9076 -296
rect 8844 -501 9076 -496
rect 7924 -962 8072 -957
rect 7924 -1056 7934 -962
rect 8062 -1056 8072 -962
rect 7924 -1061 8072 -1056
rect 7126 -1506 7252 -1501
rect 7126 -1600 7136 -1506
rect 7242 -1600 7252 -1506
rect 7126 -1605 7252 -1600
rect 2644 -2856 2870 -2851
rect 2644 -2952 2654 -2856
rect 2860 -2952 2870 -2856
rect 2644 -2957 2870 -2952
rect 7366 -3194 7690 -3189
rect 7366 -3322 7376 -3194
rect 7680 -3322 7690 -3194
rect 7366 -3327 7690 -3322
rect 2648 -3764 2874 -3759
rect 2648 -3872 2658 -3764
rect 2864 -3872 2874 -3764
rect 2648 -3877 2874 -3872
rect 12142 -3910 12296 -3905
rect 7362 -4104 7694 -4099
rect 7362 -4236 7372 -4104
rect 7684 -4236 7694 -4104
rect 12142 -4174 12152 -3910
rect 12286 -4174 12296 -3910
rect 12142 -4179 12296 -4174
rect 7362 -4241 7694 -4236
rect 12146 -4336 12296 -4331
rect 2540 -4352 2702 -4347
rect 2540 -4456 2550 -4352
rect 2692 -4456 2702 -4352
rect 2540 -4461 2702 -4456
rect 12146 -4452 12156 -4336
rect 12286 -4452 12296 -4336
rect 12146 -4457 12296 -4452
rect 7344 -4688 7716 -4683
rect 1997 -4808 2207 -4803
rect 1997 -5008 2002 -4808
rect 2390 -5008 2396 -4808
rect 7344 -4824 7354 -4688
rect 7706 -4824 7716 -4688
rect 7344 -4829 7716 -4824
rect 1997 -5013 2207 -5008
<< via3 >>
rect 5736 6198 5930 6370
rect 9558 6202 9754 6398
rect 5322 5020 5494 5190
rect 9944 5106 10040 5188
rect 2594 3716 2922 3908
rect 4844 3874 5018 4082
rect 6638 3866 6830 4084
rect 8416 3878 8610 4056
rect 10338 3898 10586 4046
rect 12048 4018 12382 4172
rect 11842 3634 11952 3724
rect 2994 3086 3168 3294
rect 1246 110 1276 310
rect 1276 110 1446 310
rect 7122 136 7248 224
rect 6906 -274 7038 -204
rect 6254 -470 6412 -286
rect 7154 -398 7254 -302
rect 8854 -496 9066 -296
rect 7934 -1056 8062 -962
rect 7136 -1600 7242 -1506
rect 2654 -2952 2860 -2856
rect 7376 -3322 7680 -3194
rect 2658 -3872 2864 -3764
rect 7372 -4236 7684 -4104
rect 12152 -4174 12286 -3910
rect 2550 -4456 2692 -4352
rect 12156 -4452 12286 -4336
rect 2190 -5008 2202 -4808
rect 2202 -5008 2390 -4808
rect 7354 -4824 7706 -4688
<< metal4 >>
rect 2592 6398 12380 6460
rect 2592 6370 9558 6398
rect 2592 6198 5736 6370
rect 5930 6202 9558 6370
rect 9754 6202 12380 6398
rect 5930 6198 12380 6202
rect 2592 6132 12380 6198
rect 2592 4486 2920 6132
rect 1558 4158 2920 4486
rect 5264 5190 5564 5238
rect 5264 5020 5322 5190
rect 5494 5020 5564 5190
rect 5264 4172 5564 5020
rect 9900 5188 10200 5346
rect 9900 5106 9944 5188
rect 10040 5106 10200 5188
rect 9900 4172 10200 5106
rect 12052 4173 12380 6132
rect 12047 4172 12383 4173
rect 1558 448 1886 4158
rect 2592 3909 2920 4158
rect 3320 4084 11452 4172
rect 3320 4082 6638 4084
rect 2592 3908 2923 3909
rect 2592 3742 2594 3908
rect 2593 3716 2594 3742
rect 2922 3716 2923 3908
rect 2593 3715 2923 3716
rect 3320 3874 4844 4082
rect 5018 3874 6638 4082
rect 3320 3872 6638 3874
rect 3320 3366 3620 3872
rect 6637 3866 6638 3872
rect 6830 4056 11452 4084
rect 6830 3878 8416 4056
rect 8610 4046 11452 4056
rect 8610 3898 10338 4046
rect 10586 3898 11452 4046
rect 12047 4018 12048 4172
rect 12382 4018 12383 4172
rect 12047 4017 12383 4018
rect 8610 3882 11452 3898
rect 8610 3878 11958 3882
rect 6830 3872 11958 3878
rect 6830 3866 6831 3872
rect 6637 3865 6831 3866
rect 3070 3295 3620 3366
rect 2993 3294 3620 3295
rect 2993 3086 2994 3294
rect 3168 3086 3620 3294
rect 2993 3085 3620 3086
rect 3070 3066 3620 3085
rect 11152 3724 11958 3872
rect 11152 3634 11842 3724
rect 11952 3634 11958 3724
rect 11152 3582 11958 3634
rect 1245 310 1447 311
rect 1558 310 8162 448
rect 1245 110 1246 310
rect 1446 224 8162 310
rect 1446 136 7122 224
rect 7248 136 8162 224
rect 1446 120 8162 136
rect 1446 110 1784 120
rect 1245 109 1447 110
rect 6218 -286 6518 -174
rect 6218 -470 6254 -286
rect 6412 -288 6518 -286
rect 6902 -204 7102 -198
rect 6902 -274 6906 -204
rect 7038 -274 7102 -204
rect 6902 -288 7102 -274
rect 6412 -290 6832 -288
rect 6902 -290 7266 -288
rect 6412 -302 7266 -290
rect 6412 -398 7154 -302
rect 7254 -398 7266 -302
rect 6412 -470 7266 -398
rect 6218 -492 7266 -470
rect 6218 -1416 6518 -492
rect 7834 -962 8162 120
rect 11152 -260 11452 3582
rect 7834 -1056 7934 -962
rect 8062 -1056 8162 -962
rect 7834 -1172 8162 -1056
rect 8658 -296 11452 -260
rect 8658 -496 8854 -296
rect 9066 -496 11452 -296
rect 8658 -560 11452 -496
rect 8658 -1416 8958 -560
rect 6218 -1506 8958 -1416
rect 6218 -1600 7136 -1506
rect 7242 -1600 8958 -1506
rect 6218 -1716 8958 -1600
rect 2524 -2855 2824 -2662
rect 2524 -2856 2861 -2855
rect 2524 -2952 2654 -2856
rect 2860 -2952 2861 -2856
rect 2524 -2953 2861 -2952
rect 2524 -3763 2824 -2953
rect 7322 -3193 7622 -2942
rect 7322 -3194 7681 -3193
rect 7322 -3322 7376 -3194
rect 7680 -3322 7681 -3194
rect 7322 -3323 7681 -3322
rect 2524 -3764 2865 -3763
rect 2524 -3872 2658 -3764
rect 2864 -3872 2865 -3764
rect 2524 -3873 2865 -3872
rect 7322 -3810 7622 -3323
rect 11010 -3810 11310 -560
rect 2524 -4352 2824 -3873
rect 2524 -4456 2550 -4352
rect 2692 -4456 2824 -4352
rect 2524 -4708 2824 -4456
rect 7322 -3910 12364 -3810
rect 7322 -4104 12152 -3910
rect 7322 -4236 7372 -4104
rect 7684 -4110 12152 -4104
rect 7684 -4236 7685 -4110
rect 7322 -4237 7685 -4236
rect 12064 -4174 12152 -4110
rect 12286 -4174 12364 -3910
rect 7322 -4687 7622 -4237
rect 12064 -4336 12364 -4174
rect 12064 -4452 12156 -4336
rect 12286 -4452 12364 -4336
rect 12064 -4646 12364 -4452
rect 7322 -4688 7707 -4687
rect 7322 -4708 7354 -4688
rect 2189 -4808 2391 -4807
rect 2524 -4808 7354 -4708
rect 2189 -5008 2190 -4808
rect 2390 -4824 7354 -4808
rect 7706 -4824 7707 -4688
rect 2390 -4825 7707 -4824
rect 2390 -5008 7622 -4825
rect 2189 -5009 2391 -5008
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1716650609
transform 1 0 6972 0 1 -108
box -183 -183 183 183
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform 1 0 7314 0 1 -352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1704896540
transform 1 0 7314 0 1 -1552
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7482 0 1 -352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1704896540
transform 1 0 7482 0 1 -1552
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_NXKS9S  XM1
timestamp 1716495612
transform 0 1 4910 -1 0 -404
box -396 -1210 396 1210
use sky130_fd_pr__nfet_01v8_NXKS9S  XM2
timestamp 1716495612
transform 0 1 10330 -1 0 -404
box -396 -1210 396 1210
use sky130_fd_pr__nfet_01v8_NXKS9S  XM3
timestamp 1716495612
transform 1 0 4932 0 1 2650
box -396 -1210 396 1210
use sky130_fd_pr__nfet_01v8_NXKS9S  XM4
timestamp 1716495612
transform 1 0 6724 0 1 2650
box -396 -1210 396 1210
use sky130_fd_pr__nfet_01v8_WWWVRA  XM5
timestamp 1716495612
transform 0 1 2756 -1 0 -3363
box -1083 -710 1083 710
use sky130_fd_pr__nfet_01v8_X7BG72  XM6
timestamp 1716495612
transform 0 1 7620 -1 0 -3717
box -1083 -1210 1083 1210
use sky130_fd_pr__nfet_01v8_NXKS9S  XM7
timestamp 1716495612
transform 1 0 8516 0 1 2650
box -396 -1210 396 1210
use sky130_fd_pr__nfet_01v8_NXKS9S  XM8
timestamp 1716495612
transform 1 0 10484 0 1 2666
box -396 -1210 396 1210
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR1
timestamp 1716495612
transform 1 0 5819 0 1 5451
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR2
timestamp 1716495612
transform 1 0 9655 0 1 5451
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR3
timestamp 1716495612
transform 1 0 2761 0 1 1056
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR4
timestamp 1716495612
transform 1 0 12217 0 1 2296
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR5
timestamp 1716495612
transform 1 0 12217 0 1 -2854
box -201 -1582 201 1582
<< labels >>
flabel space 5792 1752 6754 1948 0 FreeSans 1600 0 0 0 V2L
flabel metal1 9346 -106 9638 1884 0 FreeSans 1600 0 0 0 V2R
flabel metal1 3300 -546 3500 -346 0 FreeSans 256 0 0 0 RF_P
port 5 nsew
flabel metal1 5680 -2098 9601 -1900 0 FreeSans 1600 0 0 0 V1
flabel metal1 6389 269 6855 619 0 FreeSans 1600 0 0 0 LO_N
flabel metal1 8306 -1050 8474 1240 0 FreeSans 1600 0 0 0 LO_P
flabel metal1 12150 -1894 12300 1294 0 FreeSans 1600 0 0 0 RF_N
flabel metal1 3725 -4177 3867 -1805 0 FreeSans 1600 0 0 0 BIAS0
flabel metal1 7164 5044 7364 5244 0 FreeSans 256 0 0 0 IFOUT_P
port 4 nsew
flabel metal1 8238 5044 8438 5244 0 FreeSans 256 0 0 0 IFOUT_N
port 3 nsew
flabel metal1 720 110 920 310 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1594 -5008 1794 -4808 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 6536 -216 6736 -16 0 FreeSans 256 0 0 0 LOIN
port 2 nsew
<< end >>
