magic
tech sky130A
magscale 1 2
timestamp 1715647744
<< pwell >>
rect -235 -651 235 651
<< psubdiff >>
rect -199 581 -103 615
rect 103 581 199 615
rect -199 519 -165 581
rect 165 519 199 581
rect -199 -581 -165 -519
rect 165 -581 199 -519
rect -199 -615 -103 -581
rect 103 -615 199 -581
<< psubdiffcont >>
rect -103 581 103 615
rect -199 -519 -165 519
rect 165 -519 199 519
rect -103 -615 103 -581
<< xpolycontact >>
rect -69 53 69 485
rect -69 -485 69 -53
<< ppolyres >>
rect -69 -53 69 53
<< locali >>
rect -199 581 -103 615
rect 103 581 199 615
rect -199 519 -165 581
rect 165 519 199 581
rect -199 -581 -165 -519
rect 165 -581 199 -519
rect -199 -615 -103 -581
rect 103 -615 199 -581
<< viali >>
rect -53 70 53 467
rect -53 -467 53 -70
<< metal1 >>
rect -59 467 59 479
rect -59 70 -53 467
rect 53 70 59 467
rect -59 58 59 70
rect -59 -70 59 -58
rect -59 -467 -53 -70
rect 53 -467 59 -70
rect -59 -479 59 -467
<< properties >>
string FIXED_BBOX -182 -598 182 598
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.69 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 884.495 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
